H    �ww@                 �ww	@�iX��@                        �)B �G@H                    x   ��8Iy�8�g�8f��8�;9m+99i�`9陼9�F�9*@�9 ��9��9	��9Z:N�:+(:I�:�[:���9���9��9�@�9E�9���9��`9�&99EC98�8~f�8�x�8x   x   0v�8#��8mc�8�	9�'9�?J9K:r9�ю9�I�9���9In�9���9��9A8�9�� :� :�6�9���97��9/m�9���9�J�9�Ҏ9m9r9PBJ9�'9��	9�_�8���8�z�8x   x   Da�8`�8(C9��9�<9[`9X��9���9ϳ�9���9�7�9F��9=��9���9>h�9w��9%��9���9�9�9H��9���9F��9���9xW`9��<9� 9�F9Zb�8Y�8?��8x   x   M��8�	9��9�89�lW9V�z9�Y�9|�9�+�9��9���97��9Cp�9�9���9rq�9���9���9J�9�,�9��9(X�9��z9HiW989L�9��	9���87��8���8x   x   �49�'9��<9�jW9hqv9�=�93 �9��9�P�9���9��9}�9�J�9�g�9�L�9�9~�9<��9[Q�9��9� �9�<�9�qv9�mW9ݬ<9 '9�59�f9i#
9km9x   x   �"999J9�U`9�z9(=�9�9�9���9�ɼ9V��9��9˔�9+�9���9���9�
�9`��90�9���9Pʼ9d��9�;�9�<�9@�z9@T`9�5J9�99ac-9�s'9n'9�_-9x   x   ��`9�1r9݃9cW�9��9���9�B�9�S�95�9��9��9��9z��9��9D�90��9�9�R�9SD�9c��9%�99X�9�܃9J5r9��`9�)T9�pL9�I9�uL96*T9x   x   ॆ9�̎9���9��9��9�ȼ9MS�9��9�9m��9F��9���9���9$��9���9<�9�9�R�9
ȼ9��9��9���9̎9£�9�Y�9$<x9q�s9�s9h:x9�Y�9x   x   �?�9PD�9Y��9�(�9�N�9���9��9�~�9���9���9L��9a�9���9s��9z��9�}�9��9��9�O�90)�9���9�D�9A�9��9媔9qK�9�{�9�I�9\��9i��9x   x   �8�9u~�9 ��9D�9j��9b�9h��93��9���95 �9_2�91�9C �9��9���9���9���9���9d�9��9�9�7�9��9��9�9�'�9�*�9��9��9 �9x   x   H��9h�9 3�9-��9��9���9&�9U��9���9�2�9J�9�2�9+��9���9��9��9��9���95�9�g�9a��9|�9�-�9�h�9\�9D��9��9�g�9�/�9�{�9x   x   X��9��9���9��9��9P�9��9J��9�9�1�9,3�9;�9���9��9)
�9��9���9��9��9>��9Rq�9x��9��9W��9�x�9�y�9e��9.��9��9�p�9x   x   ���9K��9
��9�m�9�I�9{��9��9���9��9��9E��9L��9U��9���99K�9Io�9��9���9���9Y��9���9�n :T:W':��:�%::�o :���9���9x   x   �V:	3�9��9.��9g�9��95 �9��9���91��9��9? �9���9/f�9���9_��9�2�9�V:e�:��:�z:u�:7�:�:�:��:)�:�y:��::x   x   8�:a� :�e�9���9M�9R�9��9���9u��9���9a�9x�9�L�9���9�g�9�� :Q�:�:"�:JG:�1:�:�!:�j":�!:�:�1:qI:Ѿ:�:x   x   �%:^� :���9zq�9p�9ԗ�9d��9��9���9c��9�9�9�q�9Z��9�� :�$:V=:��:9:$:��):V.:�)0:�)0:].:��):v$:B9:;�:=:x   x   \�:v4�9Ύ�9��9��9��9,�9��9��9l�9r�9ڊ�9���96�9z�:�=:�y:T� :��):a�1:u�7:r;:��<:gr;:��7:_�1:~�):]� :�y:�=:x   x   XZ:���9i��9���9���9*��9�W�9_X�9���9���9���9{��9��9�X:�:�:� :��+:{5:��=:fxC:��F:�F:�xC:X�=:_{5:��+:�� :��::x   x   ���9���9�;�9��9�U�9�ϼ9.J�9Zμ9PV�9!�9�;�9���91��9Q:��:';:�):�{5:��?:�G:�L:�YN:ݥL:'�G:��?:�{5:ʷ):�::�:�:x   x   ���9�n�97��9�0�9� �9V��9���9�!�9�0�9���9�o�9��9��9��:�J:�$:��1:/�=:ȡG:5�N:BuR:|vR:��N:x�G:��=:�1:�$:�K:��:μ�9x   x   $��9.��9R��9v�9J&�9XB�9X%�9z�9���9���9@��9@z�9���9E:6:��):��7:�zC:��L:vR:RtT:CvR:F�L:*zC:��7:}�):�5:J}:���9&|�9x   x   �B�9�M�9���9}]�9C�9�C�9�_�9���9�M�9�@�9��9���9�s :v�:�:�.:�u;:ȇF:�[N:
xR:�vR:f[N:�F:�v;:9.:�:͛:�u :9��9���9x   x   �G�9�֎9}�98�z9�~v9��z9��9�Ԏ9vJ�9�)�9j8�9��9�:��:Z�!:�.0:��<:��F:ڨL:��N:��L:��F:��<:%.0:t�!:��:�:L��9;�9�)�9x   x   ���9MAr98a`9�tW9�zW9#c`9�Er9Ƭ�9⽘9A#�9�s�9���9N-:�:�p":O/0:Hw;:}C:��G:�G:�{C:�w;:�.0:�p":�:
.:���9�s�9!�9���9x   x   ��`96JJ9s�<9�$89��<9�DJ9<�`9$c�9洔9�'�9��9���9�:�:�!:.:�7:��=:��?:k�=:��7:v.:�!:":��:���9K�9�'�9뵔9bb�9x   x   �,99N'9�	9:9�!'9.99A:T9INx9wU�9�2�9� �9+��9�+:��:�:[�):j�1:�5:15:ω1:o�):�:��:O.:���9���9$5�9V�9�Ix9<T9x   x   aH9I�	9O9��	9�A9#q-9��L9�s9v��9O5�9i�9S��9!:4�:�7:� $:D�):��+:�):�!$:�7:՜:W:��9-�9�4�9���9��s9��L93o-9x   x   x�8k�8q�8��8�q9ʀ'9��I9��s90S�9-(�9�r�9���9[u :>:�N:*>:�� :d� :�=:�M:�~:sv :���9�s�9'�9sU�9��s9��I9�~'9n9x   x   Ll�8���8We�8�83-
9)z'9\�L9�Ix9��93!�9�9�9^��9��9��:��:~�:}:{�:+�:�:j��9���9�:�9  �9���9:Gx9��L9I}'9�4
9i�8x   x   �{�8���8���8���8�u9�i-9o6T9�`�95��9~(�9���9)z�9��9U:�:@:�@:2::=��9_|�9��9S(�9���98`�9�7T9�k-9zk9���8���8x   x   8Q�7!��7�u8�1q8��8�9t39��g9.A�9�@�9{|�9�o�9��9�8:�
:5]:�
:�;:���9;p�9�z�9�?�9�?�9��g9�39+�9���8f?q8@v8���7x   x   "��7g�8�JI8�k�8y(�8��9�lH9cP|9X-�9!�9�c�9���9���9{f:C�:A�:�d:P��9���9}d�93�9�-�9�R|9�hH9[�9�%�8�a�8iEI8�81��7x   x   vf8=CI8�e�8���85R	9K�39��b9�n�92��9-�9_r�9�\�9���9��9���9���9���9Q`�9�q�9�+�9ݵ�9kn�9��b9=�39�R	9���8m�8GI8�`858x   x   q8�c�8��8�:9U�)9�S9`�9�o�9>��9ۉ�92��9�3�9��9!��9��9��9?0�9���9���9��9,q�9�ހ9&�S9��)9=:9���8�Y�8�#q8.�O8��O8x   x   ۷8��8GN	9e�)9*
O9�Vx9��9���9S��9��9���9
��9���9�7�9���9���9���9���9���9���93�9�Ux9�	O9M�)9�L	9I%�8w�8���8	��8B��8x   x   �9��9��39r�S9�Tx9ʪ�9_ף9���9��9�D�9�E�9�q�9��9��9�o�9aG�9�A�9*�9藷9`գ9���9�Tx9��S9�39��9��9QI�8��8�
�8�E�8x   x   j39�bH9�b9�ހ9���9�֣9"�9�L�9�#�9�x�9
��9���9$�9���9���9�u�9>(�9�K�9��9�֣9�ߑ9�߀9*�b9�dH9�399V#9��9w�9��9T#9x   x   ��g9�D|9cj�9Kl�9���9e��9 L�9m4�9q4�9���9�2�9��9��9�0�9���9�5�9�0�9oK�9ؔ�96��9�k�9?j�9<E|9b�g9�.X9H�M9�CH9�BH9{�M9�.X9x   x   29�9�&�9��9y��9¶�9Z
�9#�9L4�9چ�9�t�9�e�9��9�f�9�s�9k��9K3�9�(�9b	�9���9���9ر�9�&�9i:�95�9O0�9�4�9�0�93�9�2�9�3�9x   x   �7�9��9{'�9߅�9o��9&C�9x�9���9�t�99��9K��9K��9���9u�9���9�v�9�=�9X��9,��9'�9��9�6�9��9c�9��9U�9-X�98��9�9��9x   x   Is�9\�9�l�9<��9_��9�D�9���9�2�9�e�9���96��9���9�d�92�9��9AG�9���9��9�m�9s[�9%t�9��9b��9���9���9oZ�9I��9���9���9���9x   x   �f�9,��9$W�9A0�9��92q�9��9��9��9C��9K��9��9��9k��9�o�9��9�,�9�Y�9���9-f�9��9Q�9���9��9���9n��9#�9i��9[O�9N�9x   x   �{�9���9���9��9h��9�9,%�9��9�h�97��9Cf�9��9�#�9��9S��9��9B��9���9]}�9+�9c�:�:�4:J�:$:-�:�3:�:��:�)�9x   x   @4:Xc:
��9��9�7�9��9���9~3�9pv�9�w�9S4�9%��9}�97�9J��9���9c:�5:r�	:�y:�:�:):+�:�:�:�:R:�y:�	:x   x   +�
:��:���94��9P��9�q�9���9p��9C��9Z��9c��9�r�9f��9r��9���9��:��
:'@:�\:�X:��%:��*:��-:_�.:R�-:�*:�%:�Z:�Z:�@:x   x   Z:Q�:���9I�9���9�J�9z�98:�9%8�9J{�9�K�9��9�9��9K�:�Y:#:�:m(:'�0:s?8:��=:�l@:�l@:a�=:�@8:��0:x(:�:�":x   x   ��
:�c:l��9�1�9���9F�9�-�9a6�9�.�9�C�9l��9@2�9���9e:^�
:�#:E� :��,:�7:��A:��I:�N:&|P:j�N:��I:�A:0�7:�,:�� :�#:x   x   ::x��9�a�9¸�9��9��9�Q�91R�9g�9k��9��9G`�9��9�8:uB:��:��,:�b::��F:'xQ:�Y:��\:��\:�Y:*yQ:��F:�a::p�,:�:xB:x   x   8��9W��9Ut�9��9s��9_��9%��9���9���9Z��9�u�9���9#��9�	:�_:(:��7:��F:wT:�V^:��d:�g:��d:�W^:JT:a�F:{�7:e(:�^:J�	:x   x   kp�9�f�99/�9Lï9ŧ9�ܣ9�ޣ9�Ƨ9�ï9U0�9�d�9�o�9�4�9H~:]:��0:��A:<zQ:�W^:,�g:�Jl:FKl:~g:LX^:�{Q:��A:�0:^:\�:�2�9x   x   |�9r�9���97w�9O�9���9��9 u�9���9�9�~�9��9�::#�%:D8:��I:�Y:��d:�Kl:8�n:�Kl:o�d:DY:��I:8E8:��%:<:��:/�9x   x   YB�9�1�9�s�9��9�dx9�ex9B�96t�9I1�9�A�9���9k]�9D :�:��*:%�=:�N:��\:�g:HMl:�Ll:�g:'�\:��N:�=:�*:w:f":�[�9���9x   x   \C�9�[|9��b9	�S9jO9x�S9t�b9'Z|9�E�9��9>�9#��9�;:#:��-:Is@:܁P:��\:��d:Ѐg:0�d:��\:��P:r@:��-:O:�9:t��9��9j��9x   x   �g9UrH93�39��)9>�)9��39-xH9��g9�@�9-�9r�9	-�9:��:��.:�s@:��N:
Y:�[^:�[^:�	Y:��N:�r@:�.:I�:P�:�.�9��9��9�@�9x   x   Z#39��9i^	9�G9\	9�9v"39FDX9K<�9'��9Ĕ�9���9�:Ş:��-:��=:S�I:�~Q:�!T:jQ:B�I:��=:��-:��:�:���9���9��9�>�94DX9x   x   T�9�7�8���8N��8<C�8��9zi#9�M9�@�9<b�9�h�9���9��:y:��*:�G8:��A:4G:�G:)�A:�G8:��*:1:��:��9Tj�9�d�9�@�9��M9Zg#9x   x   ��8�q�8i��8Uq�8]��8�i�8`�9�XH9�<�9e�9F��9�1�9b;:C:_�%:��0:P�7:�f::��7:C�0:�%:�:w::./�9Y��9Ed�9>:�9�ZH9/�9�f�8x   x   �Rq8h`I8�iI8<Nq88�5�8��9�VH9E>�9���9��9`��9�":d:pa:�(:z�,:�,:�(:�`:�:G#:���9U�95��9�?�9�YH9F�9/�8���8x   x   ߃8.�8k}8�P8�Ș8�%�8y�9ذM9�<�9~�9��9\�9�:�:�`:q�:8� :��:Ya:#�:q�:\�9��9u�9"=�9U�M9��9,�8֘8KP8x   x   ꨻7Ӳ�7O)8�	P8u��8?]�89b#9�>X9 =�9��9���9{�95�9o�	:�E:3':)':E:�	:d4�9V�9���9q��9->�9�>X9(b#9^�8l��8�P8p-8x   x   di~�ki���)��[���7��8A2�8�999�|9�O�9rs�9�	�9�*�9|z	:,:�A:W:q}	:�+�9O
�9�q�9�M�9��|9;99�3�8B��8q:�7H��E�)��i�x   x   �i�4�?���ٷ�}c6MM/8q�8�
9 �R9i��9��9u��9&�9�=�9#�:��:��:��:
9�9��9���9��9ۼ�9��R969`x�8�V/8��a6c�ٷ��?�oi�x   x   U�)���ٷ4��L� 8!��8Df�8��59��q9jB�9���97��9_��9�/�9t�:�}:�:3�9¬�9z��9��9}C�9�q9��59�g�8J}�8�� 8��w�ٷZ�)��=�x   x   .���_ib6r� 8�Ǌ8|�8m%9��[9@u�9S��9���9�2�9N�9�8�9��9��9�9�9D��9=1�9���9׈�9�u�9i�[9�%9�|�8�̊8�� 8e�`6o��J'Ϸq<Ϸx   x   �ʥ73/8s|�8�w�8��9JkQ9$�9���91�9�B�9���9D��9��9T2�9Z�9���9m��92B�9��9���9|�9�kQ9"�9Oz�8�t�8�D/8��7_\�6���5���6x   x   �y�8B_�8QY�89�$9ZiQ9ऀ9PA�9��9�&�9��9��9r@�9��9C�96>�9`�9;
�9%�9ڂ�9h@�97��9�jQ9��$9�[�8�b�8�m�8e�G8�2$8]#$8��G8x   x   ��8Z�9�59��[9a�9�@�9f��90H�9S��90i�9��9���9H :���9���9�e�9���93G�9��9[A�9��9��[9C�59�9��8ی�8S�8خ8��8��8x   x   .)99��R9O�q9�q�9��9�~�9�G�9���9bF�9t��9���9?�:��:8��9���9�F�9���9AH�97�9��9�p�9��q9�R9L(99��%9�]9'�9�96`9��%9x   x   i�|9ŵ�9�<�9��9q�9�$�9���9DF�9�}�9���9H�:�:! :L��9`}�9RE�9���9�$�9�9���9=�9˵�9��|9�k9�O^9��V9X'T9��V9�P^9�k9x   x   �E�9\�92��9��9�?�9I
�9�h�9}��9ٛ�9:b:`G:YF:�b:���9��9�h�9"�9�B�9���9��9?�9�D�9�f�9�r�977�9T��9}��9�7�9�q�9�f�9x   x   zh�9���9���9e.�9���9��9���9���9��:�G::�G:��:���97��9h�9���9,�9N��9ҵ�9�i�9׾�9v`�90�9�f�9}6�9�c�9L�9b�9���9x   x   T��9b��9��9]��9F��9�?�9���9��:t:G:H:�:U�:���9?�9���9���9~��9���9���9'��9T��9���9Ep�9�^�9U`�9�r�9*��9x��9Ą�9x   x   ��9k5�9;*�9�5�9��9�9�H :��:d:�c:u :��:vG :P�9+�9q8�9�,�9�1�9��9{�:}�:�:s�
:a:� :`:��
::�:Z�:x   x   Ku	:i�:)�:��9d2�9�9���9���9���9/��9���9���9��9p2�9k�9��:h�:yw	:S�:��:N�:W�:LP#:�J%:\K%:eP#:֟:��:�:c�:x   x   � :��:�{:��9��96A�9���9x��91��9���9e��9�B�9��9��9,}:��:��:7:�!:@�):�1:�8:�<:�p=:�<:�8:��1:U�):�!:�7:x   x   +>:Y�:F�:�:�9���9��9k�9�L�9nK�9�n�9��9h��9v<�9�:��:O>::T�(:��4:ҿ?:�I:3�O:�NS:�MS:��O:�I:#�?:\�4:�(:�:x   x   |:o�:$3�9� �9���9�9���9���9���9j�9���9�9=2�9��:]::ix+:_S::șH:�0U:Z
_:]Le:�rg:�Me:U	_:'0U:K�H:�T::w+:�:x   x   �{	:68�9���935�9�G�9!,�9O�9�P�9X-�9uK�9u4�9���99�9�z	:�9:i�(:�T::��K:�y[:�h:/r:�w:<w:�r:��h:Iz[:�K:�S::r�(:�9:x   x   *�9��9���9���9��9��9ȯ9���9��9���9N��9�	�9B(�9��:z!:�4:*�H:�z[:��k:��x:Zn�:ց:�n�:��x:��k:�{[:�H:y�4:�!::�:x   x   �
�9n��9�9x��9���9�I�96K�9���9���9N��9T��9W
�9H�:o�:x�):c�?:;4U:��h:�x:M �:7�:h�:��:��x:�h:�2U:��?:/�):H�:��:x   x   �s�9��9�I�9N}�9L�9��98�9�{�9I�9��9�v�9���9M�:�:Q�1:�I:W_:r:�o�:��:ڳ�:��:p�:�r:�_:�I:R�1:^�:n�:���9x   x   �P�9	9��q9�\9>~Q9NQ9"\9��q9�93R�9PͿ9�	�9L:!�:08:/�O:�Re:�w:�ׁ:��:��:�ׁ:�w:�Re:;�O:�8:d�:�:
�9#ο9x   x   ��|9W�R9�59�%9/�9�%90�59��R9��|9>u�9-p�9���9�
:�X#:O<:�VS:�yg:Pw:0q�:t!�:&q�:�w:T{g:�US:�<:�X#:�
:���9m�9�x�9x   x   ZD99Q9���8&��8+��8ą�8�9�A99�3k9Q��9�!�9��9Pj:T%:�y=:�VS:�Ue:�r:g�x:��x:�r:WTe:dVS:�y=:�S%:�j:H��9�&�9��9~.k9x   x   ZF�8Ώ�8���8h�8���8틹8�E�8_�%94l^9	G�9-x�9fq�98
:U%:�<:��O:�_:ıh:\�k:j�h:�_:K�O:�<:WT%:�	:Kq�9�r�90G�9r^9m�%9x   x   ���8-�/8�8�8v�/8���8���8
w9R�V9=��9�G�9�r�9�i:-Z#:J8:�I:K8U:L�[:|�[:l7U:�I:�8:�Y#:ok:tq�9}L�9k��9p�V9�t9{��8x   x   Mv�7<Cd6w
��d6u�7ZH8y�8��9+CT9��9�t�9ۄ�9#�
:Q�:��1:��?:�H:��K:8�H:��?:�1:�:��
:���9�r�9��9�DT9n�9D �8?H8x   x   I��]�ٷl�ٷ[��2�6�w$8u �8m�9q�V9�F�9}"�9f��9�:��:��):"�4:z[::�Y::��4:k�):r�::,��9i&�9-F�9Y�V9 �9X��8Qs$8�9�6x   x   ��)��}?���)���η!�5�`$8��8�u9i^9p�9Zq�9'
�9�:��:!:��(:�|+:	�(:+!:��:��:�
�9:l�9?~�9�m^9�p9��8�k$8.��5D�ηx   x   ��h�#�h�,�=�>�ηU?�6�H8E��8��%9:,k9�r�9�ɿ9g��90�:��:�=:$:B:�<:[�:��:��9�̿9jv�9$(k9��%9ܨ�8��G8��6��η��=�x   x   ö ���������ոs��.�4�MU8��8OpO9(�9.Ⱥ9T�9�� :C�:��:qY:	�:��:�� :��9�Ǻ9a|�9]pO9] �8oU8��4������ո'�����x   x   ���F��Pj�8�����uG�7�D�8;9ORl9��9��9E	�9���9�:�}:H~:ɇ:)��9	�9��9{��9*Sl9<9�>�8�c�7"��7����k�-�����x   x   8���n��=��:�F�!C5��p8D��8F9W�9��9@��9�U�9���9z:zC:V:i��9�W�9��9��9��9]F9к�8{�p87<=5t�F�U3���l�Q�����x   x   ��ո�����F��=���<?8(��8]).9]�r9��9��9��9!��9I��9\:�:���9���95�9��9��9��r9i+.9���8h??8m�����F�ç� �ո�N�BS�x   x   f'��=���>5�3?8���8��"9�b9Mi�9Q�9�l�9s4�9fS�9�� :��:� :�S�95�9Ck�9�P�9i�9m�b9��"9��8E0?8�895�����������6����x   x   �t5����7��p8g��8��"9�]9�ڌ9s��9�5�9~�9��9)��9K:�~:���9��9 �95�9���9=ی9C�]9�"9���8�p8��7��5����Ur-��x-���x   x   ��T8�+�8���8�".9F�b9�ٌ9e��9�\�9y��9�&�9��9%�:Z:*�:ߴ�9�$�9���9�[�9��9�ڌ9�b9s$.9���8 '�8��T8��7�h7!7��h7L��7x   x   ���8,9�F9<}r9�f�9�9j\�9���9c�9y :P�:�: �:9�:e :�b�9��9^�9~�9�g�9d~r9�F9{,9���8�\�8%	�8Q�8�T�8��8�]�8x   x   �ZO9Al9�x�9i�9)N�9 4�9��9	c�9W" :��:�
:�:��
:Z�:." :b�9���9
5�9^M�9��9x�9hCl9�YO9�~89F0(9�l9�+9�f9j/(9V�89x   x   s�9d�9��9��9�i�9�|�9�&�9� :�:AW:��:��:
W:��:v :c(�9{�9~j�9�99�9L�9�q�9o�9��9�]{9NEw9�Kw9�_{9��9�n�9x   x   ;��9Q��9��9��9�1�9��9e��9��:��
:=�:4�:J�:Y�
:O�:��9��92�9N�9ށ�9���9��9݆�9N�9��9���9���9���9.�9��9w��9x   x   � �9��9�N�9���9�Q�9D��9ܷ:�:�:��:��::��:��:���9�P�9���9�O�9* �9%�9:��9���9��9�@�9k4�9\5�9�@�9���9��9!��9x   x   [� :��9���9���9^� :�:X[:��:9�
:�X:z�
:��:�Y:�:�� :��9��9���9�� :��:lW:��
:7�:��:�S:P�:��:F�
:�U:�:x   x   �:��:��:e:\�:b�:2�:��:��:�:$�:�:��:v�::��:-�:�:j�:b�:�L!:T':1Y+:�-:ם-:�W+:+':�L!:c�:��:x   x   ��:�y:�A:�:L� :���9x��9{ :K% :e :4��9��9� :�:B:.z:R�:w*:r�):d�3: =:yQD:�	I:��J:�I:(RD:c�<:��3:w�):m*:x   x   U:�{:� :7��9X�9��9�+�9�j�9�i�9�/�9�9sV�9���9N :0{:�U:	%:�2:��@:��M:&�X:P�`:m�d:}�d:��`:��X:��M:��@::�2:�%:x   x   ��:S�:���9J��9;�9���9(��9 ��9ۤ�9��9u:�9���9դ�9�:w�:=
%:�#6:��G:=�X:7tg:s:lz:��|:Bmz:�s:�sg:��X:%�G:�"6:�
%:x   x   s�:���9fZ�9�$�9�r�9>�9�e�9yh�9�?�9�t�9�$�9�Y�9���9)�:�-:��2:�G:SD\:�o:v�~:��:}χ:χ:r�:�~:�o:�C\:��G:��2:�-:x   x   � :�
�9Ѝ�9	��9�Y�9��95��9���92Y�9��9��9�9l� :��:L�):��@:�X:%o:qL�:H�:q��:�U�:���:,�:�L�:^o:�X:��@:�):��:x   x   ~�9Q�9@�9O!�9/s�9��9��9�t�9�!�9���9�
�9J�9��:7�:��3:,�M:�xg:��~:�:|��:�C�:C�:n��:%�:��~:xg:��M:��3:a�:��:x   x   �ʺ9��9|��9��r9X�b9[�]9��b9��r9F��9R�9�˺9���9�_: U!:�=:*�X:s:��:��:hD�:�,�:rD�:��:��:\s:��X:x=:XS!:�^:���9x   x   ǀ�9s`l9�+F9�?.9��"9��"9 ?.9r-F9bl9��9a��9	�9��
:�':�ZD:��`:nsz:�҇:	X�:�D�:(E�:�W�:|҇:fsz:u�`:�YD:�':��
:)
�9d��9x   x   ){O9�J9���8"�8!-�8�#�8��8J9zO9���9H)�9,��9��:�c+:�I:��d:D }:�҇:���:���:h��:Ӈ:� }:��d:@I:�b+:��:&��9'�9]��9x   x   �7�8�\�8Gq8�?8Ê?8�Iq8�]�8'5�8\�89/��9�9	V�9�:;�-:��J:��d:�vz:|�:s�:��:��:duz:p�d:��J:/�-:�:�V�9��91��9՛89x   x   �5U8�֟7ZFN5�3��a�N5�̟7�<U8���8dR(9��{9^�9�J�9\_:��-:!I:S�`:qs:��~:@P�:�~: s:��`:I:��-:�_:>I�9x�9w�{9�U(9��8x   x   �J4��d�V�F�\�F��b�]R4�l��7�D�8�9kw9�Į9�K�9��:�c+:�]D:W�X:}}g:�o:4o:A}g:O�X:�[D:0d+:��:eI�9�Ȯ9vlw9	�9tD�8_��7x   x   �����������������L��j7���8�L9qw9�9�V�9R�:�':`
=:	�M:ȧX:�K\:+�X:\�M:�=:�':��:[W�9 �9�kw9�O9⌚8�vj7�M�x   x   ��ո<Y�V�C�ո�ԣ�Z$-�Ȓ7ۊ�8 �91�{9��9D��9��
:rW!:��3:?�@:G�G:J�G:��@:��3:�U!:#�
:���9��9��{9W�9i��8|�7�"-��ѣ�x   x   w��C��+���7�V��&3-��*j7DE�8L(9�9�)�9�
�9q_:��:I�):*�2:�)6:8�2:�):�:`:z
�9�%�9��9_P(9J:�8�7j7�+-����9�x   x   C��������@��أ� [��g�7x��8��89�|�9���9Z��9>�:��:�1:�%:�%:p1:��:��:���9Z��9��9��89��8���7�g��ڣ��=����x   x   �J������>x���V�<�'��ԸP���f5X8a�9�7w92I�9ɇ�9u1 :�":�:��:�:�!:31 :(��9J�9�4w9y�9(JX8 ��w�Ը͜'���V�k=x����x   x   !����~���c�h�;�$��ꇸ�7�H�8[r:9�S�9V�9.��9��9|�
:��:g�:s�
:��9}��9�R�9�T�9Gx:9�B�8T}70ㇸb���;�^�c���~�v��x   x   wCx���c�H�A�n,��W��k����^p8J�9ZGg9��9���9�S�9V��9��:�
:��:���9wQ�9���9��9XAg9S�9ip8|���Wc���-���A���c�uCx�!�x   x   @�V��;��.��"��G���0#8���8��H9(��9�E�9E&�9Ț�9D�:�:O:��:��9.'�9;D�9���9�H9ە�8	#8����j��!.���;�S�V��d��d�x   x   Z�'��$�Na��Q���[1
8d��8R89r��9�Q�9)_�9Z9�9�9�m:��:�m:��9�7�9^�9ZR�9#��9oK89���8 A
8���m���!��'�f<��	C�9<�x   x   ��Ըe���֓�K#8��8V39��|9쫢9\t�9/*�9��9ps:V�	:�	:ns:��9�,�9^v�9Z��9-�|9s39���8��"83������� �Ը��4�� �����x   x   Yo����7�7p8���8SN89?�|93�9a�9��9;M�9�G:KM:eW:�M:�G:�M�9��9;�9��9��|9�G89ڄ�8�>p8�7����kEx�R����>�������Nx�x   x   �W8w(�8.�9��H9��9ê�9�9z�9^�9�':��:�^:�]:��:�':�^�9~�9��9���9i��9N�H9��9� �8~�W8��7���5y��}���ޒ5P�7x   x   ��9^_:9/9g9`��9�N�9!s�9h�9?^�9�:�:f:��:�:d�:��:]]�9�9�t�9�P�9s��93g9�c:9 �9��8���8+ק8���8>Ч8���8`�8x   x   ]w9YI�9���9�@�9�\�9G)�9M�9'(:f�:o:�E:YE:�:}�:�(:O�9�+�9[�9�?�9+ �9J�9iw9�^9�yK9�7?9d9999�8?9�sK9^^9x   x   �:�9K�9���9!�967�9��9\H:��:=:SF:"�:kF:�:�:/G:��9x4�9[#�90��9PI�9�:�9#ʣ9;˝9`Ù9e��9��9G�9wř9W̝9�ȣ9x   x   =y�9$��9;L�9���9��9�s:�N:;`:O�:�F:G:�:�_:�O:�s:-�9 ��9:K�9-��9�z�9q��9��9}w�9��9�'�9�'�9���9tv�9���9���9x   x   V* :���9���9��:�m:��	:gY:S`:�:�:m:�`:�X:%�	:�m:��:���9���9* : $:[�:��:W

:��:�A:��:�

:��:N�:�$:x   x   ^:��
:�:M:q�:2�	:�P:$�:��:O�:c�:�Q: �	:��:>:�:ʬ
:!:��:�9:L�!:+"':�?+:�m-:*l-:h>+:F"':��!:19:��:x   x   0�:�:d�
:�:�o:�v:�K:�+:��:�,:`J:�v:�o:D:��
:��:��:�":��,:6�6:CJ@:��G:�L:�5N:��L:��G:�I@:�6:��,:�":x   x   q�:�:F�:t�:�%�9�"�9JW�9Xh�9g�95X�9;$�9]%�9y�:(�:ҍ:�:��(:rv7:EF:��S:�6_:y�g:��k:��k:�g:6_:d�S:yF:w7:L�(:x   x   �:^�
:L��9B��9�?�9t6�9��9n��9e�9{6�9�>�9���9���99�
:+�:�(:�2;:P�M:!`:.�o:DT|:l�:fw�:��:�U|:��o:l`:��M:K3;:��(:x   x    :���9�U�9�.�9h�9 ��9��9��9���9�g�9�/�9�V�9��9�:� ":]y7:��M:#>d:
�x:���:dɊ:z�:�:�Ȋ:u��:E�x:3?d:��M:�x7:� ":x   x   �0 :���9��9�M�9�]�9S��9���9 ��9�^�9HN�9��9Z��9�0 :��:W�,:�F:n`:͗x:k��:�I�:N��:*Z�:��:wI�:/��:]�x:�`:�F:��,:��:x   x   M��9uX�9P�9�	�9��9B
}9
}9�	�9=�9Z�9�Y�9U��9`,:�A:y�6:�S:9�o:h��:�J�:�Ζ:��:p��:�Ζ:iJ�:��:��o:ҿS:1�6:�A:U,:x   x   |N�9#\�9=Ug9<�H9�f89�239�f89��H9(Ug9�[�9xM�9���9��:��!:#S@:�>_:[|:̊:��:���:�ߜ:���:]��:�ˊ:�[|:�>_:S@:z�!:�:��9x   x   �@w9��:9�9���8�.�8�/�8���8h�9+�:9@w9�ޣ9Н�9��:�,':��G: �g:� �:��:�\�:��:ü�:R\�:��:� �:��g:��G:�-':��:��9Lݣ9x   x   ��9�g�8O�p8�n#8�
8?t#89�p8hf�8%�9 7^9G�9���9@
:�K+:��L:��k:+|�:�:6��:�Ж:Ð�:w�:�{�:��k:-�L:�J+:�
:4��9�9�6^9x   x   ͅX8��7�ْ����0��N˒��7��X8+]�8]�K9�ڙ9���9D�:<z-:&BN:B�k:"�:Z͊:M�:M�:�͊:�!�:��k:GAN:fy-:K�:���9�ؙ9��K9<a�8x   x   ��������q:���鼸�:����;����7�7�F�8�c?9-��9A�9�N:Ly-:c�L:��g:�`|::��:���:�_|:,�g:p�L:�y-:$O:�?�9X��9�c?92E�8q0�7x   x   x�Ը}
��|�W
�{�Ը^�w��5S%�8�699�ϖ9�@�9 �:�K+:A�G:�A_:w�o:Z�x:��x:+�o:�B_:,�G: L+:��:�?�9Ж9799�'�8f��5�w�x   x   �'�(�;��A�d�;�A�'��|����ʺ��C�87999a��9O��9a
:�.':�U@:��S:S`:�Gd:r`:��S:IV@:h/':c
:���9���9�599kA�8����à�,}�x   x   s�V���c���c���V�6
<����U�������8p`?91ۙ9r��9[�:;�!:�6:�F:PN:�N:F:��6:��!:��:��9�י9�_?9K �8p��������h<�x   x   /8x�Ѵ~�d9x�L�d���B�	��aʠ�'��5;�8.�K9��9���9��:hC:@�,:�7:g:;:~7:��,:�C:�:~��9���9�K9�6�8$_�5�͠�4��`�B�U�d�x   x   �������~��d��<�w����w�Oϴ7"R�83-^9ڣ9|��9�-:��:u#":�):�):�$":��:-:���9ڣ9�-^9�K�8Wٴ7��w�*���<��d���~�x   x   ]U˹��ǹ�3������5{]��k	�x	 ��u�8p�19W9Æ�9R%�9��:'\:�:\:��:�$�9��91ď9��19�q�80��o	�iy]�?�����1����ǹx   x   ��ǹO[���y���ۚ��)y�]�-�����V]7#j�8in`9���9�c�9���9��:��:G�:��:���9�e�9N��9l`9�x�8 ]7�����-��)y�=ٚ�Uy���]��/�ǹx   x   ;6���z��n�������A�f��5F��r�8�J39h��9�O�9���9g�9�t:�
:Lt:�e�9���9�P�9��9�C39f�8?'������A�������oz��5��)��x   x   ��"ޚ����?H�j���7�+?V8�i9�v9���9zn�9���9c�:�	:3�	:��:R��9�q�9ͅ�9��v9'l9�EV8��|���RH���<ܚ�/���8���6��x   x   �����0y���A������
5�)U*8c97Kd9���9���9
<�94=:�p
:<;:gp
: =:�8�9d��9W��9�Nd9.9�N*8:�4�����v�A�k1y�]���xf������&h��x   x   @�]�&�-���฀��M*8�V9�n\9kU�9u�9F{�9B:�l:�:�:�m:B:�|�9Px�9\R�9�l\9�\9_M*8�*�����-���]���}��@���?��� ~�x   x   ^|	��4������X'V8<9|m\9��9_��9p��9�:R�:E:��:AE:	�:�:��9���9C�9�k\9�9�+V8N}��A6��p�	���/��sG�7dO�rG���/�x   x   sY �i]\7��8)b9Gd9�T�9H��9U��9��:(�:�!:d�:��:":��:��:���9���9nR�9�Id9�f9��8�\7{I ��ϣ�p�ܸE�������I�ܸ�֣�x   x   �G�88F�8�=39Ŋv9���9ht�9���9��:��:CN:P�":�C%:j�":0O:�:��:u��9�u�9���9�v9�839/N�8�H�8���7E����lŷ����1Mŷ�^�����7x   x   "�19[`9���9h��9���9P{�9:��:�N:�o$:��(:ױ(:�n$:O:��:�:��9v��9��9���9�[`9D�19�94@�8���8��8qؠ8鑴8�:�8I�9x   x   
��9��9�H�9�j�9;�9�B:��:#:��":m�(:��*:��(:��":�":n�:B:Y7�9dn�9CH�92~�9Ҵ�9�5�9�@h94-W9�M9b�I9M9�.W9�Ah9|6�9x   x   oy�9Z�9��9���9c=:8n:'G:��:�E%:��(:p�(:�E%:��:>G:�n:+>:X��9���9eZ�9�z�9m�9�9'��9�f�9S�9-ߦ9Qd�9ť�9��9�k�9x   x   ��9��9\b�9��:�q
:(�:��:��:��":�q$:� #:��:��:[�:q
:W�:�_�9Y��9��9W��9]��9��9RJ�9	��9�\�9a��9�K�9���9j��9���9x   x   $�:�:Fs:g�	:X=:p�:QI:q&:NS:�R:w%:AI:l�:�>:��	:Et:n�:��:)
:�>:<�:w:��:::a�:�:,�:�=:d
:x   x   �W:��:��
:ڪ	:�s
:er:)�:�:1�:3�:Y�:�q::s
:ߩ	:�
:
�:�W:X�:� :��':C�.:?�4:�B8:C�9:lB8:W�4:I�.:��':: :$�:x   x   ��:?�:du:��:�A:�G:":4�:��:t:G:uB:��:�v:Z�:��:�X :w,:e8:݄C:�1M:A<T:��W:��W:�;T:@1M:؅C:8:0,:�X :x   x   QZ:_�:�j�9���9�C�9���9?��9��9\��9���9�C�9\��9ri�9W�:�Z:FZ :0:�@:X�P:)�^:��i:��p:�hs:K�p:��i:l�^:3�P:֘@:;0:�Z :x   x   ��:���9X��9\|�9���9F��9���9���9S��9���9�|�9~��9���9U�:��:�	,:��@:�U:��g:�w:-f�:�T�:[T�:�e�:�w:��g:�U:>�@:�,:S�:x   x   `'�90l�9�Z�9���9`�9�b�9T!�9�c�9��9��9�X�9�j�9�&�9&
:� :O#8:ΝP:��g:�G|:�:��:�Ȍ:��:��:�H|:<�g:��P:$8:� :A
:x   x   \��9*��9��9q�v9>od9y�\9��\9�nd9R�v9O�9���9l��9q��93G:��':��C:l�^:��w:��:�]�:!)�:7(�:�]�:��:Ùw:��^:w�C:;�':cE:��9x   x   �ˏ9[�`9K^39-�9979�9�59�9�`397�`9�ɏ9	��9#��9K�:��.:V:M:��i:�h�:��:�)�:�>�:�)�: �:�h�:	�i:.:M:N�.:��:��9\��9x   x   �	29���8�=�8��V8��*8
�*8��V8>�8��8�29vL�9!��9��9�:��4:FT:��p:TX�:}ˌ:�)�:�*�:ˌ:2X�:� q:FT:��4:4:���9:��9�K�9x   x   ��8�^7	E�����_s4�!���P����^7"��8d�9cph9ٽ�9bc�9\�:XN8:m�W:4rs:\X�:��:`�:P�:�X�:mqs:��W:�M8:A�:ve�9z��9_vh9T�9x   x   ���쩸q�����8���ێ��쩸e�����7���8�^W9m��9M�9:ȗ9:U�W:�q:�i�:	�:3�:}j�:�q:e�W:��9:_:��9�~�99XW9���8��7x   x   �\	���-��A�!�G�)�A��-�?]	�)���MX�����8�9M9v��9}w�9K:-O8:TGT:N�i:��w:�O|:��w:��i:HT:�N8:�:�w�9���9�AM9�8Bͻ�:���x   x   Ni]��y�%������>y��f]���/�;�ܸ"ķ�;�8f�I9���9��9p�:ՙ4:�<M:��^:R�g:��g:c�^:X=M:y�4:�:��98��9��I9o7�8O�÷ޫܸ��/�x   x   �됹Tњ�����Қ��됹j�}�[UG��w���\��,/�8�;M9�|�9�d�9:��.:q�C:d�P:JU:[�P:d�C:��.:):_e�9�}�9�>M9:3�8nk��n}��tVG���}�x   x   ��Ds��Bs���	���\���4���HO�΁���+ķC�8ZW9a��9���9Q�:&�':�&8:��@:^�@:w(8:��':��:F��9f��92RW9s�8�"ķY����CO��5��\��x   x   �.��5Y���/��>2��⍡��5��ZG���ܸ�U��&��8Ehh9}��9P��9G:�# :�,:: 0:�,:s" :dF:��9&��93mh9|��8�����ܸ�\G�u7��x����1��x   x   /�ǹ��ǹa���1���a��n�}�p�/�;������7�9�F�9�|�96��9
:޺:X^ :�^ :��:�
:d��9-}�9�E�9�9{��7Q���y�/���}�m_��t3�����x   x   ���[�	��?��o����ٹ�L�����#+��n�VHa8q0*9���9�Ӷ9�z�9:@�9��9�A�9u�9:Ҷ9��9�6*95Na8�n��!+����I����ٹ�q��?�M�	�x   x   �	�ǵ��)���X⹢�����J�L�����$�7�9��m9���9�t�9���9�(�9�'�9y��9w�9��9��m9�
92�79���һL�g��H���	T��(�������	�x   x   �@��*��&��Rƹ�䞹�a�X���X�84T9��9�R�9��9��9L� :���9:��9�M�9��9�:T9@�8������(a�>㞹1ƹ 幊*��K@��{�x   x   �r���Z�ƹG���9j������˷!�8O�D9ݕ9�9y��95� :z":�$:�� :L��9)!�9�ڕ9$�D9��8i�˷����9j��H��ƹ�U�ts��E�����x   x   ��ٹR���枹%;j��	����r�8��<9M��9��9���9�:G�:,:f�:(:��9)��9a��9ǆ<9��8Z��r�	��;j��䞹4���e�ٹ� ��x   x   �Q�����Va����G����8�.99���9 r�9:��9��:n�:"�:-�:X�:Ɖ:݀�9�s�99��9�,99|�8z��_��7a�x ���L���ʹ��ԹB�Թʹx   x   �Ȉ���L�t��̷��8�.99Z��9rD�9���9*�:R:�J#:�X&:�J#:.O:��:���9VE�9�Ñ9 ,99i�8�	̷��+�L��Ɉ�JU������d��:��kQ��x   x   :1+������u���8��<90��9�D�9d��9�:}<:��):��/:�/:��):}<:��:+��9�B�92��9��<9q�8���t���I.+���e��醹�1���3���솹��e�x   x   mBn�Ю�7�8ϳD9y��9s�9��9��:7�:UE-:��5:��8:��5:_F-:1�:��:���9�s�9%��9A�D9w�8���7xVn�K��QG(���D��N���D�\I(�y��x   x   	a8W9�.T9~ܕ9��9���9��:�=:"F-:��7:ԋ=:3�=:S�7:F-:�>:��:��9���9<ܕ9�0T9�9�a8��ʶ1r]�8��?�Ը8�Ը�@���a]��z˶x   x   !*9E�m9$�9��9]��9��:ST:B�):��5:ٌ=:)@:�=:	�5:�):nT:�:@��9<!�9\�9Y�m9N#*9��8Ԉ~8Vu�7c^�6�u�����6�h�7��~8��8x   x   ���9���9RR�9Ŕ�9��:v�:3N#:g�/:��8:g�=:�=:��8:J�/:�M#:��:��:Y��9�N�9���9���9��`9�;69ȳ9�"�8�f�8�c�8J�8S�9�;69��`9x   x   �Ͷ9�r�9E��9]� :��:N�:�]&:$�/:��5:�8:j�5:~�/:�^&:E�:U�:/� :���9�u�9�ʶ9�96��9���9Q�x9��m9;�i9`�m9��x9v��9���9��9x   x   �v�9���9���9�%:�0:��:�P#:z�):�K-:�J-:��):P#:��:*2:�&:���9M��9Dt�9���9���9[�9���9�Z�9.��9N°9UY�9��9���9��9���9x   x   �>�9v+�9h� :R):J�:�:?V:�C:��:UD:/Y:n�:��:�':)� :-+�9@�9�)�9=��9���9�j�9]��9���9���9ͦ�9a��9�j�9"��9c��9	)�9x   x   O��9--�9���9�� :R�:��:��:�:��:z�:��:��:� :���9�-�9��9�u�9j��9�:�:��
:"�:�,:�,:�:��
:
:+:��9w�9x   x   �E�9���9��9��9Ҷ�9ђ�9��98��9���9���9[��9���9��9���9�E�9�x�9r:;:PZ:��:� :}�$:u5&:0�$:�� :O�:�[:m::s:7x�9x   x   4|�9���9\�92�9��9���9=Y�9DV�9B��9=��9r1�9S]�9���9R�9s2�9���9�<:��:-I#:�%-:�D4:��7:c�7:�C4:�'-:_H#:��:P=:D��9)4�9x   x   ܶ9u��9��9T�9��9A�9�ؑ9��97�9t�9��9���9�ڶ9���9��9x:�]:�J#:U1:qD<:�9C::�E:m:C:C<:�T1:�J#:�\:�:?��9���9x   x   �ĉ9�m9�^T9��D9�<9NX99�W99�<9��D9�YT9+�m9�Ɖ9�9��94��9:}�:�(-:�E<:�G:'�L:޺L:�G:�E<:P)-:��::���99��98�9x   x   'R*9�+9}c�8�U�8�l�8bj�8�l�8�\�8�d�8S09N*97�`9G��9/�9�{�9K�
: � :I4:y<C:��L: P:e�L:�;C:dI4:�� :��
:Z{�9�	�9���9��`9x   x   [�a8�%�7��^�ʷ$���b�ʷ�����7��a8�/�8�g69�˅95��9���9��:��$:O8:(�E:R�L:}�L:�E:�8:
�$:��:1��9,��9�ǅ9�f69�4�8x   x   C�m�h���B�񸬸��	���ΐ�_���U�m�v,ŶO?8��9�y9[p�93��9�5:>=&:�8:?C:�G:�=C:F8:3<&:&6:���9�q�9� y9��9�A8��Ŷx   x   +���L��`��j��j���`�y�L�+�Ǘ��\����7�8��m9]ְ9��9�5:3�$:oJ4:�G<:CI<:UK4:��$:\6:��9pذ9Y�m9Ip�8���71�\���x   x   ����}��Ԟ��8��7Ԟ� ��|���ve��(��ⱸ���6���8"*j9ذ95��9<�:U� :.-:zY1:V,-:m� :Y�:{��9�װ9�)j9%��8�$�6�汸�!(�Lye�x   x   &?������`�Ź^�Ź����k=���D��M؆��D�2]Ը�;�����8��m9�m�9a��9A�
:X�:�M#:�N#:��:��
:��9p�9��m9��8�ݻ�(hԸV�D��Ն��C��x   x   ��ٹ�J⹰�乞J�:�ٹAʹ���"���N��~Ը�}�6�b�8$y9O��9+{�9B:Ta:ޓ:[_::�z�9İ�9�y99a�8�Y�6�oԸ{�N��$�����{ʹx   x   l���!���"���j��-����ԹaX��)&��_�D�:���r�7
�9�ą9@�9���9�:�>:�?:�:c��9A�9M9��9^�7����h�D�'���S��x�Թ:��x   x   _=�\���=����k�m�Թ ��Tᆹn0(���\���~8WW69���9���9!��96��9Fu:^��9<��9}��9��9�U69��~8��\��1(�;܆�E	����Թ���x   x   ��	�Q�	�&z�[�����'ʹjI��u�e�n��O�ȶ\	�8��`9��9���9�.�9.z�9Kx�901�9���9��9:�`9��8��ȶ�����e�FL���
ʹE�蹐��az�x   x   UR6� �4�][/�R%&�Z������o�b��������z �m�g�8�8���849�C[9��h9�F[9�49���8q�8��g�>| �����ā���n湂�����&&�5[/��4�x   x   ��4�n0�I�'�p���D	��蹕P��b)��z��Ȉ��}8	�9
�d9eP�9|��9��9tR�9�d9!�9��}8K��ŝ��*��3N���蹔E	�g����'�Ln0��4�x   x   \/���'�D*�i�	��E蹂嵹r}�������Y]�8�@9Ύ�9�۪9��9M��9��9�ڪ9�9�	@9�a�8�x������}�w嵹	B�k�	�e-���'�#[/�M�1�x   x   �%&����O�	���㱴�Y�v��.��*�.��"�8��b9'R�9>��9bv�9�X�9�\�9�w�9��96T�9��b9�8�91�A(����v������{�	�C��>'&���+� �+�x   x   ���yD	�E�L���Jdt���.�7�09B9L��9���94!:��:	:�: :'��9��9�9�69M7U��jdt�豴��A蹴F	���	�"�>�%�X�"�x   x   "�����㵹I�v�в�=g7�9��9О�9��9 &:J�:�#:�#:+�:�&:T��9S��9m߈9�9��f7.��i�v�䵹;蹚�� ��h������x   x   o湫N���|�W#��*7�9\5�9�*�9~� :�R:%(:�+3:��6:`+3:�|(:jS:� :�,�9�5�9�9Z�7 "����|�uO��n湑��	��������Q��x   x   ׀��^&������n,��89�9�,�9(�:+:�X0:Gx>:��E:��E:ey>:EY0:�:�:�+�9��9�696�-����#��\���F�G����c��d�v���R�x   x   ����u��f���:�8 9��9�� :I:�3:�]D:�$O:��R:�#O:=^D:�3::8� :i��9�9�:�8�/��������������Jٹx�﹅�������Mٹ����x   x   Br ��W�{�8��b9���9��9�U:,[0:�^D:gR:۵Y:��Y:,fR:�^D:�[0:GU: ��9��9��b93z�8]j��p ��x���.���0˹ڹ�ڹ42˹�*��|��x   x   �g���}8 @9�\�9���97+:��(:|>:�'O:V�Y:�_]:W�Y:B(O:|>:j�(:�*:���9�^�9�@9��}8ug�r&�4���A��Y_���k��YY���C��5���&�x   x   �8�9���92��9�':��:�13:��E:��R:��Y:ٸY:�R:,�E:H13:$�:�':Ʋ�9�9ȼ9�8z͍�$��<n��ɐ�k杹�杹s͐�w;n�m$�ȍ�x   x   `#�8��d9��9��9ϋ:�#:�6:_�E:n)O:�jR:I+O:��E:��6:-#:
�:p��9��9�d9��8��j7Q��������Q���t��[�� �t���Q�]��X���nk7x   x   }349Z_�9��9k�9�:>#:\43:��>:\eD:�dD:~�>:-43:�#:L:�l�9��9�^�9`249��8k�����[���>-�}�A��A��C-�5��3ߔ�+�i���8x   x   �`[9Ù9��9�q�9��:�:�(:�b0:X3:�b0:�(:V:͍:oo�9b��9|Ù9Gc[9�9��g8�%��J���qԸ�W����AV��kԸ`S��B��+h8 9x   x   [�h93ř9[�9)��9�,:�2:�^:o$:c%:f]:�1:-:n��9:�9ƙ9&�h9�=!9�̾82r8��<��3E�I/������œ��D.���(E��<�uv8ӻ�8�>!9x   x   n[9i�9��9���9D�9��9� :G�:d� :���9$�9���9$��9f�9\m[9�B!9.�8|�t8V�7���$����5�K�H�a5�£����F�7 �t8P9�8?!9x   x   �?49:�d9^��9�o�9���96��9pF�9�C�9��9a��9�o�9a��9~�d9�E49R(9J߾8y�t8��85'P7PO���h�|Ť�Ǣ��8�h��nM��)P7��8��t8�־8�+9x   x   �N�8�99A@9l�b9yH9��9�O�9���9�I91�b9C@9��9�N�83!�8�.h8Ȧ8�I�7�cP7V�6 ��5�;�p�8�Q#����5#�6�P7<:�7��8g>h8/#�8x   x   9�8"i~8/Ҷ8���8�o9R9�P9�g92��8Ͷ8{c~85�8��l7�Q����%�;�1��zM�g
�5��6���6��6�ɒ6[��5v2N������;�C
�4iZ��m7x   x   :�f����ͻ��#��7SJj7*�7��!��̠���� �f�����Y[��1ǔ������D�T!��I~h��;����6��7���6@��FIh�v��o�D��"�������Y��'���x   x   �L ��j�W��޼���L�R����ɺ�cj��I �I�%���#�ӂ�P��EԸZ����4�����f�7�1��6ڻ�6��6�c`���4����I7Ըb��?����#���%�x   x   Q������0�|�"�v��3t�Μv���|��������f��&#��n��wQ��&-�;C�3o��Q�H�Ut��V)�	��6���un��A�H�Sk��L�+%-��oQ��n��$���h��x   x   �m���8��fϵ�雴�r����ϵ�<��n���鴹����2������S�t���A�g���z��=�4�L�h�1��5/��5�h�]5��q�����A���t������4��W���괹x   x   �]�f��!/�>蹒/���繪]����<ٹ:#˹�R���ڝ��Q����A��I���V���N�M��T�6KP��k��>���S���A�S��ٝ�	N��\#˹�<ٹB�x   x   ���)>	���	���	�]?	������������dڹb��Tޝ��t�U9-�>^Ը�E�WA���O7��O7����<E�VԸ�2-�4�t��۝�f���ڹ/���������x   x   ���ˤ��'����|�����$���^�'���hڹ�R��Ȑ���Q���2T����<�¹�7��8���7J=��O�������Q�Ȑ�T��
ڹ�|���`�>��V��x   x   <#&���'���'�%#&��"����N���a�{��.˹b@���7n����攸�a��C8�xt8�ut8RC8����딸���I4n��@���,˹���b�ɑ�Ɇ� �"�x   x   FY/��k0��X/�5�+���%������j����Kٹu)��55���$�崙��t��g8H��8�8x��8�g8M/~�i���:$��5��T*��NIٹ���E��<����%�i�+�x   x   F�4�Ǡ4���1�~�+��"���������u����}��"&�|ۍ�N4j7Ｉ8�9d#!9�!99ҩ89hj7)ꍸ�&��|������A�|�������"���+��1�x   x   a�e�Lmd�U^`���Y�[>P�_�D�[�6��9'������.�5	͹�^��ګ��}/��x���|/�����wa��~	͹K�B��H��_9'���6���D�>AP� �Y��^`�Cmd�x   x   imd��&`��W��~K���;�$�)��<�$m����ӹ� ��µ����>���"?���藸�闸<����0�>�շ���!���ӹ�p��<�9�)���;��{K�s�W�s&`��nd�x   x   �]`���W���I��&7��� ����۹X����a�,������M8�-�8ۇ�8o�9?��8%�8a�8��6���8�a��W���	۹���"� �i'7�i�I���W��\`�rAc�x   x   <�Y��|K��%7�N��`� �83ù�z���	��'��k��8+^290�z9T��9�f�98g�9���9�z9�\29���87����	�&y���7ùG� �����$7�zK���Y��`���`�x   x   =;P�6�;�� ��� ��κ���b�PQ���e8^�79�?�9Ź�9_��98��9���9���9���9ʹ�9�>�9+�79�e8R���b��˺�^� �@� �>�;�C<P���\�a���\�x   x   @�D���)�����+ù��b���u��;�8�u9�\�9ـ�9g:�e:�&:�&:zf:ef:���9�]�9��u9�>�8��u��b��,ùb����)��D�TBW���`��`��BW�x   x   ,�6�5���ڹ�n��V.��FN�8t��9���9��	:X$:m8:�<D:�\H:?<D:�8:-X$:T�	:M��9���9VS�8�#���n����ڹ�5���6���O��_�e�I�_���O�x   x   W0'��Y���E����	�re8��u9���9U3:�"/:^�G:��X:�a:�a:��X:Z�G:n#/:g3:���9;�u9�de8D�	��F���Y��z0'��F�AF]�U�h���h�pF]�9�F�x   x   P����ӹŐa�cٞ�89�j�9Z�	:P%/:'KM:�xc:�q:.�u:�q:�xc:�JM:�%/:_�	:�k�9�	89�➷*�a���ӹ���؞<�rpY��pk�؅q�ok��qY�O�<�x   x   �������H���8�U�9R��9_$:��G:�zc:HFv:��:�:�Ev:�{c:~�G:H_$:z��9
S�9w�80G��������E?1��8T���l�LVy�Yy���l�}7T��?1�x   x   R�깞�����g�29���9Cr:x8:��X:q:�:�_�:�:�q:��X:�8:r:���9�29��ȗ�����Z%�]�M��}l����" ��ӫ�w~l��M��Z%�x   x   ��̹�:>��87{9S��9�r:�GD:��a:��u:2�:�:��u: �a:�GD:�r:���9y7{978�6>���̹���9�F�bk��H��4و��و��I��8k�h�F����x   x   �7�����1Ȱ8���9���9�#&:�iH:��a:q:�Kv:�q:�a:>jH:�#&:"��9���9/Ͱ8=��8��V&�t�?���h��������	��4���t���	�h�η?�%�x   x   ��������l-�80��9?��9�%&:JD:��X:O�c:�c:C�X:�JD:>%&:���9I��9�&�8o���G����e��E9�`f��$��i�&���}��� �S$���f��F9�2g�x   x   ���H5��NE9-��9v��9x:8:~�G:^UM:�G:�8:iw:���9Đ�9�H9�6�����J ��.4� �c���1���7������w7����/����c��,4�? �x   x   �͎�/��L>�8iɖ9A��9�x:�h$:a1/:�1/:�h$:^y:���9&Ȗ98�8
/��ώ�&�����0�N�a�����xG��C����;���;������>G�������a���0�����x   x   ����}��{�8�R{9���9���9#�	:�A:_�	:��9m��9*O{9��8�|��������B�/�S�`����/6��w��#[������\�����K6������`���/�����x   x   �|��T��Pr8��29�h�9̃�9���9���9܃�9�f�9�29no8����|��� �a�0�O�`����4��4���rt��������vs��>����3��>����`�+�0�� �x   x   ]2��t!>��^��`�8�389dv9P��9v9�889.\�8�c�@ >�#0��Gc��-4�C�a�Z���]4��1���;��q�º��ź�º���*���!4�����Y�a�,4�d�x   x   (�̹,���K������Vf8���8���8b6f8���� ��?�����̹;#�vD9��c�6���7��'������gĺ��ɺ�ɺ�eĺR�������6��g���w�c��E9�� �x   x   ��깋���fa�C�	�G���h�t�����	��ga�����7��)����?�`f�����H��I��Zv���º��ɺI;̺��ɺΪº�u������I��g���f�J�?�{��x   x   ���c�ӹX1���T��X~b���b�V��~2��2�ӹ���MW%���F�ݷh��%������ä�*^��?���ʒźN�ɺ��ɺԑźw���_���ä�?���&��S�h�!�F��V%�x   x   ��aM��J�ڹ�ù����ùh�ڹ�I�����;1��M� k�%������:���?��]�������%�ºqiĺb�ºΑ������=?��];��(������6k���M�9<1�x   x   �*'��,������ ��� ����7.�+'���<�
8T��~l�dJ������ޖ��@���2A���a��Zy��\��E���y���a���@����������!����J����l��6T�5�<�x   x   Ӯ6�ʇ)�4� ���6� ���)���6�^�F�	pY�u�l�z��7܈��������=���Ǥ�������!���I������Ȥ�7>���������?܈������l��pY���F�x   x   `�D�F�;�Y7�7��;���D�t�O�^F]�=sk��Zy��#��Dވ��Í���������KO���>��Q<��O<��>��4P������`����Í��݈�$��q\y��tk�=D]���O�x   x   �:P��tK��I��tK��8P��@W�n�_�#�h��q�I`y�H���O��<���,�����ū������ ��G�����4���,������ O����_y�o�q���h���_��@W�x   x   ̚Y��W���W�I�Y���\�Z�`��e���h�tvk���l�Q�l�-+k���h�f���c�R�a��a��	a���a���c�e f���h�q+k�V�l�a�l��yk�K�h��e���`���\�x   x   |\`�$`�[`�`�`��a���`�/�_��M]�4{Y�'CT���M�8�F�Y�?��Y9�kA4�1��/�O1��A4��Z9���?���F���M�`CT��zY�QK]�]�_���`�5a���`�x   x   {ld��md�Ac���`���\�GW�0�O��G�4�<��L1�j%����8��{��* ����5���+ ��z��6���ui%��L1�:�<�-G�7�O��FW�>�\��`�8Ac�x   x   ����~���O��%�����O��茺�ߍ��&�� ����'��6���"��`(��Zᖺ9&���ᖺ�'��/��ܫ���'��Y����%��kߍ��猺N���������O���~��x   x   )~��_Ɋ�䩇��y���X}�ZTs��i���`�@�X�Y�Q���K��?G���C��zA�
F@�sF@�{A��C��?G�	�K�.�Q���X��`���i�mUs�X}��x��񩇺�Ȋ�o~��x   x   IN��ܨ������Wo���Z��E��)1����b��������Z͹D����r��Wk���n������\͹��K��������&1�4�E��Z�/o�����ި��uN��N���x   x   0���v��$o��oR�.3��@����nү���z���$�N��x��G\&�I��74g�7[p'����M��_�$���z�6Я���� E��-3�AnR��o�\v������������x   x   ���_O}���Z��)3��	�tν�i[�L3���P8-59H8p9�j�9�9�@�9��9Tj�9�6p9�19}�P8}/���m[�n˽��	��*3��Z�CP}����Ѕ���g�����x   x   �G��MFs� �E��7�Ž�Rf.��3�7n�;9��9$�9&�:��:Nj:Zj:T�:s�:�&�9���95�;9_4�7sg.��ƽ��9���E�cEs�hG��gs��D?��O>��zs��x   x   Bތ��vi��1���EB[��҉7��i9.��9�I:�0:�$F:RpS:k�W:oS:&F:�0:�G:%��9��i9���7�C[�ı�w1��wi��ތ��L���Ԫ�a®��ժ��K��x   x   Ӎ��m`����㬯�w����;9���9�k:zYE:^d:ςx:tT�:JU�:#�x:d:LZE:�l:���9��;9Ó�+�������o`�Ӎ��Х�I���\v���u��÷���ѥ�x   x   ����rX��z�t~z���Q8�9�R:^E:;n:���:�l�:�I�:�k�:ط�:�;n:^E:�Q:Ϥ�96�Q8��z��{��qX����8����aú�Ѻ�pֺG�Ѻbú����x   x   ����0�Q�����[$���9�H�9:#0:� d:���:�ؒ:�\�:�\�:sْ:e��:pd:�#0:�I�9%�9�^$������Q�芐�Eĳ�1cкD�����@��S���bк�ó�x   x   �����K��a�}X���p9��:J5F:��x:Cp�:�^�:l�:�^�:o�:1�x:F6F:��:�p9)S���_�y�K��������/ݺO���� ����[ �����1ݺi���x   x   /����G�H͹���褖9;�:��S:�[�:�N�:�_�:�_�:�O�:O\�:Y�S:��:J��9ˮ�J͹�G���������p��-�8�����Q������,��o�y��x   x   �����C�<��֝�w.�9��:��W:�]�:�q�:~ݒ:~q�:U]�:d�W:��:Q2�9���;���C�T���?�ƺk���b�����&���)�4�&�/���������ƺx   x   ���)NA�z ��LU�7ꁯ9?�:�S:C�x:���:+��:g�x:�S: �:/~�9�5�7� ��|MA�F��2x˺�F������p(��5�.�<���<�`�5�"p(����G���x˺x   x   Dɖ��@�?��+�7�6�9�:�=F:*d:�In:�)d:P=F:=�:7�9�O�7����@�'ɖ���κ����F��22��!C�5�M�ՃQ�1�M��!C��32�:G�Q����κx   x   ��@�X��O)�ح�9v�:�-0:smE:�lE:t.0:�:���9ϗ �����@����(�к�1��� ��9��5N�,�\�kid�id���\��5N���9��� ��1�Z�кx   x   �ɖ��NA�9��\�ݻp9�_�9g_:t:�_:�]�9��p9�k��7��:MA��ɖ���к���j@#��>�9V�gh���s���w�n t�Cgh��V���>��@#�g��J�кx   x   !���C��͹W*����9ྦ9��9���9Ӿ�9C�9F%���͹q�C�����κN2��@#��*@��<Z���o�t%�����8����$��o��<Z��)@�A#�3���κx   x   �����G�X�$?$���R8�0<99Qj9�,<9(�R8B$�X��G�U���Qz˺1��m� �c�>��=Z�AKr��{���j���s���j���{���Jr��=Z��>��� ����q{˺x   x   ���"�K������\z��P����7(=�7�X���^z�q���r�K�뗓���ƺ�J���I���9��V���o�,|��������\�����4|��(�o��V�]�9�!J��J���ƺx   x   �����Q�gv�e����
[�j.�x[�핯�"v�ŇQ����&��q���9���62��9N�Ckh�.)��k��c��&���h��"l���(�kh�:N��62�����������x   x   ����oX����f��W������
��R���oX�C�������iv�A ��u(�l'C��\��t�>���?v�����D	��%v������t�F�\�.'C�Lu(�� �jv� ���x   x   ���m`�s1�)0����}-�S1�hm`���ȳ��5ݺ 2�:!�j�5�Z�M��pd�lx�Ι��n��<���m��򙃻�x��pd��M���5��!�1�M6ݺGȳ�x   x   =ԍ�Kui���E�G3��3��E��ti�5ԍ�����}iк�������&�&�<���Q�Srd��	t��-�{�����.�=	t�+rd�S�Q���<�L�&� �����iк����x   x    ߌ�iDs��Z�vbR�m�Z�hBs��ߌ�wԥ�'hú�亹&�����)���<�m�M���\��qh�9�o�Tr��o�yqh��\�4�M�t�<���)����&�9���hú�ԥ�x   x   vG���K}��o�� o�$M}�1H���O��F�����Ѻ������Э&��5�j-C�PAN��(V��GZ��GZ��(V��AN�-C�F�5��&�U�������0�Ѻj���dP��x   x   7���t��ڀ���t��9��Hv��ڪ��~���{ֺ��}(� ���&��{(��?2�"�9��>��5@��>��9�@?2�|(��&�����(����zֺT~��*ڪ��v��x   x   �������������� ����C���ɮ�����Ѻ��亢���)7���5���S�i� �JM#�=M#�7� �GT�����y7�1������4�Ѻ*���Uʮ�C��<���x   x   �N��Ȋ��N��ƥ���k��_D��Iު�ö�pú�sк"Dݺń麵���O`�����>�
�(?���C_���������:Cݺ[sк�pú�¶�bݪ�kD��Em������x   x   ;~���~��X����������{z���U���ݥ�<̬��Գ�ز���!��/�ƺ�˺��κ��к�к}�κ��˺z�ƺ�!��屺��ճ��̬�8ݥ��V���z������}�������x   x   �g��x���ބ��Ȧ��dM��E�Ǻ��պ-溈m������{�&��H� ���&�K�*��),�P�*�i�&�� ���`|�4��)m��[-溨�պ��Ǻ�M��������q���x   x   J���b���]��-���Q�����u���.����º��̺��ֺߊຖ����x��ү���̨躸����ֺj�̺��º/����$����䠩��]��֘������x   x   u����Z���C���F��j_��@���kc��~[���[��z��姍�������C���TD��ҥ��5������"�������\��g\��<b�������_��GG��EC���Z��삭�����x   x   .��������C��� ��|�z��\�F�B�K�-���V������	�2�����a������	�$����B���-�P�B��\���z�* ���C��'���z��������x   x   �B������CX����z��5I�"����޹^����8��/ø���=�6��7�t8���7��6���0øS�8��^����޹���	4I�s�z��X������EC���Ǻ5q˺��Ǻx   x    �Ǻ�����w��_�\�[���~��rn�;��8�_9���9���9J��9���9���9$��9���97��9x�_9���8�n��}��&��9�\��w��������Ǻ�#ں������$ںx   x   ��պ���S��S�B�,�޹$J��I9���9��:�!5:��M:N\:1�`:�\:��M:�!5:��:���9�L9G���޹8�B�zR��x��ުպh��/� ������ ����x   x   6�g���F��8�-�t(��D�8(
�9r�$:�|Z:��:���:Aȓ:�ɓ:���:5�:�|Z:?�$:�
�9�6�8)����-��F��V���溉����)w��v�b��
�x   x   P����º�B��I���b8��W`9�
:��Z:&��:
��:�s�:&T�:�q�:���:մ�:�Z:
:�Y`9�[8���bC����º�O����8�$�*�/���3���/�<�$�s�x   x   ����̺i犺�T�������9<95:P�:n��:���:�K�:BL�:+°:U��:��:�95:k�9�����U��抺��̺��/�!�&�8�#I��tQ��tQ�I��8�'�!�x   x   �h�>�ֺه��9����/��9� N:���:�y�:IN�:q��:>N�:�x�:Ψ�:zN:���9\�����x����ֺ<i�ܻ0�,gM�+�c��rq�]4v��rq�l�c��gM���0�x   x   ����dຜ\����4�6��9<\:>ԓ:*\�:�P�:2P�:G\�:�Փ:�;\:�9#"�6B���\���d����?�g�a��6~�!9���{���{��69��#6~���a�7?�x   x   n� �`�躥В����CF�7� :Y�`:�֓:�z�:Ȱ:�{�:�֓:R�`:1 :�r�7���В�'��d� �W#L���t�+������������:�������t��"L�x   x   /�&��f�I������n�8) :B>\:`��:ֺ�:˺�:���:x?\:c :��8Œ�!���{f�S�&�L�V����ꂗ�A���z��2h��Mh�����޺������b���v�V�x   x   y�*����J��p�����7�9lN:��:þ�:Y��:$	N:y�9ɛ�7��������񺇸*�Z�^����W���絻�ƻ�Vл��ӻ�Vл�ƻY赻B�����r�^�x   x   -,��񺄁����NB�6|��9�E5:��Z:ޖZ:&F5::��9{�6��͂��J���,�8�b�����ާ��!���.Իڅ⻅ �n 껵�⻶.Ի�!���ާ����?�b�x   x   ��*��i�Qђ�����i����9F:�$:�:n��9IN�����ђ��h�*��b�jt��m��ߝƻHD޻Z��U���+ ��U�����C޻�ƻ>m��Kt��Пb�x   x   $�&�����^��������5�`9�3�9�6�9�`9<���R���^����躩�&���^����m����Ȼ���*��������������w����㻍�Ȼ�m��i����^�x   x   u� ��h�̉��S�P:8��Ђ8!�9�Â8�58�mS�/���4iວ� �j�V���6᧻ßƻ��Ե��q(��c�����c�b(�������*�ƻ�৻���"�V�x   x   >��;�ֺg芺���j��H����������N芺��ֺ����(L�G������K%���G޻����-)�lJ����[��fJ�J)�̣��_G޻,%��@�����{(L�x   x   �m�a�̺�D��g�-�.v޹�L��u޹Z�-�|D��~�̺�m�$?���t�������3ԻT����Ne�^��æ�^��Be���a��4Ի�������t�$?�x   x   �����º�G��̤B�d��e����B�G����º���l�0��a�����j���yƻό�j\��������G������Z\���⻏ƻ�������.�a���0�x   x   `X�����SQ��ѱ\�� I���\��Q��p��XX����!�:pM�DB~�犙�?
��C_л6	�;0 ����Pg�M�g����[0 �	��^л�
������A~��pM��!�x   x   �溭	��tu��ށz���z�"v�������C�)�8�͌c�@@��)$���q����ӻ�
�`��I���,��,�t���_���
�1�ӻpq���#��A@���c���8���x   x   ԰պ����V�����fV��=���պ��ض$�vI��q�샎�����r��.bлP����&���������ʳ𻗑��aл�r��������J�q�I�T�$���x   x   ��Ǻ����A��XA�������ǺE�������/�i�Q��Dv�S���I&��_��$"ƻB;Ի?P޻w��k��UP޻U;Ի/"ƻ���S&��3���Dv���Q���/����Ũ�x   x   �G��5����@��ꜩ��G��=-ںE� �߀�f�3��Q���q��C��ŏ��KǨ�N����.��ɪƻ��Ȼ��ƻ�.������]Ǩ�ď���C��=�q�Q�Q�o�3����'� ��-ںx   x   ڣ���[���Z��뢳�n�Ǻp��m����U�/��I���c��K~�����T���^��	짻�y���y���맻�������G���L~���c�JI��/�������㺑�Ǻx   x   냭�����1�������z˺���.� �n���$�O�8�_{M���a���t�󫂻������������j��t�����t���a�e{M�7�8�Y�$������ ����|˺���x   x   u�������L������H�Ǻ?3ں��"�n%���!���0��3?��9L���V���^���b�/�b��^�* W�Q:L��3?���0���!�U%�&"�����3ں��Ǻ�������x   x   #�Ⱥ2
̺�ֺ"u�%��������f�4��K�Td�{}�A���}���x��ލ��)L��ۍ���x���}��A��}��Sd���K�Զ4�J�������0u纵�ֺ%
̺x   x   �̺��κWԺ��ܺ���n�����>��z#��3��C���R���_�q�h�+jm�3jm���h��_���R���C��3��y#�������������Z�ܺ�WԺ��κM̺x   x   |{ֺ�RԺF\Ѻ��κ�|κ@@Ѻ��׺ʺ�+��(
�rk�!)���N�݃��(�k�e
�=��+�q��&�׺D@Ѻ|κ��κ�[Ѻ^RԺ6}ֺ)4׺x   x   i���ܺ��κ�俺����%��vM������\��\V��\c���䫺4��+�����Z4��y䫺�b��W��6]��ѿ���M��D%��x����俺2�κ��ܺ�g纺 �P!�x   x   )���,��7pκj���R���w���K���*����������Φ���T�����,S���������{����7�*���K��w�tR������pκB��G����e����e�x   x   P
�0���\,Ѻ����v�5
(���ƹe,�V|ӳ�8d�H9�-u9��9i�9�0u9��H9��8��-a,��ƹ,	(���v����[,Ѻ8����	�W��ew!�hw!����x   x   ��������׺�7����K�^�ƹ�4����9S��9��*:�ZG:/2W:�+\:�1W:FXG:��*:*��9���9V6��	�ƹ�K�7����׺-��2���'3��?�~�C��?�Y'3�x   x   v�4������z���]*���+���9I�:�g:�͍:�m�:���:N��:�n�:�͍:�g:4�:5�9��+�Y]*�0��������Y�4�SO��qb�jfl�ifl��qb�@SO�x   x   ̲K��a#����S8��@q���5���9��g:���:8%�:���: }�:O��:\%�:���:�g:���9,�5�p�I8��� �ia#�H�K�W�n��܄�Ti��ZT��hi���܄�S�n�x   x   �5d��t3��� ��+�����[��8��*:�ٍ:�*�:�p�:m��:Q��:~q�:�)�:Yڍ:�*:���81��9,��;� ��t3��5d����o+�����㺭�Ⱥ�����Z+�����x   x   ��|���C�w�	��3���3����I9i�G:�}�:w��:���:�D�:���:���:�}�:7�G:q�I9�2���3��}�	��C���|��:���_���F»
�ͻ�ѻ"�ͻ�F»�_���:��x   x   �.���R��M�c���?����?v9�fW:���:���:q��:���:߈�:I��:5gW:�Bv9`���ͱ��vM�h�R��.���ک�rsƻ\޻���������c��m޻{sƻ�ک�x   x   [j���c_�6
���������~�9�c\:엦:v��:Az�:��:藦:�a\:]�9��������X
��c_�Pj��Kq(ۻ���^��F��� F�c�����^(ۻx   x   �d���h��d��鳺�c���~�9WjW:���:�3�:3�:y��:5kW:׀�9�c���鳺�d��h��d���iŻ<&���Lx�� "�ư'���'�� "�@x�
��n&�~iŻx   x   �y���Fm�K���곺'����Mv9��G:a�:��:��:ِG:HMv9���B곺u��|Fm��y���Yλ� ������$��<3�1O<�Rl?�2O<��<3���$�Ο�� ���Yλx   x   �8���Gm��e�P��^���J�I92�*:�g:5�g:I�*:��I9k���� ��f��Gm��8���ӻ� ����u/�IhA��FN�u U�~ U��FN�FhA�"u/����� ��ӻx   x   ]{���h���F����4����8�*�9� :(�9$�8�1��̴������h�v{���ӻG�����-6��K��E\�F�f���j�@�f��E\��K�26����A���ӻx   x   xg���h_�?Q�Y6������ F51J�9�M�9��F5G���6���P�bh_��g���\λE�S��i8���P��-e�i�s��c{��c{�b�s��-e���P��h8�W��N��\λx   x   7n��A�R���	�/��)j�_�+�d�����+�@j�/��z�	���R�In��,nŻ�%��N��!6���P��<h�s{z�#�����)��`{z��<h���P�"!6�C��k%��enŻx   x   �3��ͰC�R�Q:��T*��aƹcƹS*�:��L���C�_3��B���-����x/�P�K�0e��|z��䄼�䈼�䈼�䄼�|z�	0e�L�K��x/�����,�9���x   x   ��|�|3���o����K�^�'�8�K�Z����+|3�{�|��᩻�0ۻǘ���$�ymA�eJ\���s����Y刼�押W刼�����s�oJ\�pmA���$�ޘ��0ۻ�᩻x   x   k@d��h#�ǝ��5��K�v� �v��5�����]h#�p@d�OB���|ƻ
���~�WC3��MN���f�ki{�C��*戼1戼Q��li{���f��MN�yC3�`~������|ƻB��x   x   ��K������׺����G�����+�׺>����K����3i��޻6��:("�hW<��U���j�k{�X��焼C��
k{���j��U�CW<�H("�Q���޻Ui�� ��x   x   ��4���/Ѻ񮱺����/Ѻ�����4�o�n��4��wR»���>N�ҹ'��u?�R
U���f�C�s�%�z�N�z�V�s���f�P
U�v?�ι'�)N����WR»�4����n�x   x   ,��9����pκ*߿�qκ�������
`O��儻����ͻ
���Z���'��Y<��QN�=P\��7e�pEh�p7e�<P\��QN��Y<���'�l�����)�ͻ����儻`O�x   x   z����κ
�κ�����23�ށb��s���ǭ���ѻ���]P��+"�GH3��sA�L�K�C�P�B�P�b�K��sA�kH3��+"�=P������ѻ�ǭ��s�� �b��23�x   x   z���g�ܺ[ѺX�ܺ֕������?�yl�6`��Gɭ�B�ͻ���6 �ۃ��%�/�/��*6��s8��*6� �/��%�ȃ�M ���`�ͻOɭ�l`���xl�T�?�L��x   x   �q纣VԺ�UԺip��m�!�!���C�({l�Iv������X»�޻/������ի�������������ҟ�����޻�X»��v��{l���C��!��m�x   x   1�ֺ��κ9�ֺX,�Z����!��?��b�lꄻ<;���q����ƻ0>ۻP=��7��s�A�����7���<�M>ۻ��ƻ�q��J;���ꄻ�b�Ӑ?�z�!�Y���,�x   x   �
̺^	̺W;׺.�o�Y��b93��iO�s�n��(���L������,Ż{oλ7ӻӻ�oλqŻ$��\�L��r(���n��iO��93�^���o��-�;׺x   x   2X�r,�����=}�DN-�z�I���l�Ta��gݠ��踻�Dѻ!e�d���_0��3�����3�I0�W���1e��Dѻ5踻�ݠ��a����l���I�N-�5}�Z��^,��x   x   ;(���{����D{��6 �+63���J�P�f�����0ܓ�EѤ����������`˻]л�\л^`˻��������:Ѥ�1ܓ�	���_�f�I�J�63�*7 �1{� ��}��'��x   x   l�������-��P�����$�gS4��G�f�[���p�[��q򉻩 ��a�������&��q�p�4�[� G�{S4�a�$�;��dP�.���8�����t��x   x   7s�gs���ɐ�������x���3{�-��������j&�-.�Wo2��n2�C,.��j&�܀�B����z��������y��������s��r�����x   x   �>-��) ��F�p�����޺��ú������Λ��뛺s���ӥ��ª������ê��ԥ���i꛺nΛ�����F󮺈�ú�޺?����F�) �F?-���5���8���5�x   x   ��I��"3�������R�ú�ǒ��DS�o��gɹ3���I�W�N+9���.���.�p$9�	�W����jɹ����CS��ƒ�Y�úD������c#3���I���Z�o�c��c��Z�x   x   �tl�l�J�^�$�����ۮ��,S��K���K�7q]�9EZ:[�':�::�"A:�::��':�Y:c�9}/�7M��<.S�vۮ�����E�$���J��tl�Z���p��fz���o��X���x   x   HO��Qbf��64��c�����@����7��:��c:��:A}�:?��:[��:}�:��:!�c:�:�/�7ƶ������c�'64�9bf�cO�����$ū�U(���(��\ū����x   x   �Ǡ�낻��F���������ȹM��9��c:���:'��:j��:|��:4��:n��:��:M�c:.��9��ȹ ���˃�y�F��ꂻ�Ǡ�����_jϻzfܻB��Zfܻ>jϻ����x   x   Qϸ�#œ��[����~���!	��Q�:���:`��:6\�:��;��;H[�:���:���:��:
��J��������[�6œ�*ϸ�:�ڻi���+�c[
�Q[
�,�i��o�ڻx   x   t(ѻ����o�p�MZ�֟��iV�K'(:Õ�:���:�;r�;(�;���:\��:�$(:�fV�H֟��Z���p�V����(ѻ����_������&���)��&����2������x   x   fF��z�����A&�T�����7��L;:��:R��:G�;O�;j��:j��:�M;:]w7������A&����{���F軰G��$��6��|D�b�K�I�K��|D�C�6��$��G�x   x   �}������;ى�p.��|��	?-�xA:q��:M��:"h�:��:���:yA:�B-��~���.�zى�Ƹ���}�����R7��tO�*@b��1n�;Jr��1n�(@b�jtO��Q7����x   x   ��C˻<玻�D2�p���<-��R;:c��:���:���:,��:�R;:�A-��n��]D2�N玻 C˻���'�vH�w�e��N~���������k��������N~���e�tH�Ӊ'�x   x   A#��?лj���#E2����u7�0/(:��:�̪:D�:�.(:�q7�Y���VE2������?лQ#�P0�!U�Y(x��d���X������Ւ�������X���d��:(x�@!U�E0�x   x   ����@л鎻j.��bRV�F�:� d:6!d:�:/VV�B����.��莻�@л����4��l]�/����S�����9���?������Z���-����l]���4�x   x   �$�F˻/܉��E&�a؟�������9{:4�9����؟��E&�Q܉�$F˻�$�Ն4��D`��%�����	K������B�ļ��Ǽ*�ļ����
K������%���D`��4�x   x   n"��������I_�������ȹ�Q�7݄�7��ȹ촛�5_��������v"�0��n]��&��.��.����ü4-м2�ּL�ּL-м��ü'��;���&���n]�0�x   x   ����7���5�p����#��� �����������������p�]���z���O�'��%U�S������3���VƼg.ּ�I�6�㼧I�`.ּ�VƼ1��l��a����%U�H�'�x   x   �O軘����[�؇�e���S��S�}������ӛ[�l����O�D���H�/x��� N���ü�/ּ
�㼏�꼝��!�㼨/ּ֘üN��� /x��H�B��x   x   �2ѻy̓���F�f�Yծ�|���)ծ�{f�2�F��̓��2ѻN��Y7��e��i���#��ߚ���0м�L��������mL��0мݚ���#���i��D�e��Y7�N�x   x   _ٸ�5�n>4�������ú�ú�����=4�򂻏ٸ�d��%$��~O��Y~��^�����ļ_�ּg�㼉��x��m��q�ּ�ļ ��_���Y~�e~O�8$����x   x   Ҡ�Anf�\�$�e���7�޺*���z�$�of��Ѡ��ڻ���7�lLb�� �������Ŵ�%�Ǽ��ּ=O�r��MO���ּ�Ǽ�Ŵ����� ���Lb��7������ڻx   x   �X��T�J���2����������؝J��X�����z��h��T�D�7@n�����S����ƴ���ļ5м"5ּ%5ּ 5м��ļ�ƴ�E���~���3@n�J�D�U��>z�����x   x   ��l��+3��I��J��,3��l��Ý�Bzϻ6�;�&�ٗK��Zr�d���������П��9�ü�^Ƽ2�üџ��������x����Zr�ǗK�C�&�16�8zϻ�Ý�x   x   �I�51 �����[0 ��I�����aӫ��xܻ�f
���)�<�K��Cn�R��c���)���T��M ��S ���T��x)��$c��V���Cn�D�K���)��f
��xܻ�ӫ�����x   x   �I-��x���by�OJ-���Z�M|���8������g
���&�x�D��Rb��b~�5o���������"��������Bo���b~�Sb���D���&��g
�J�໫8��|����Z�x   x   �{����5��5{���5���c�3���h:���|ܻK9�F���
7�g�O���e��<x�b����/���/��q����<x���e�r�O��
7�/��a9�H|ܻ::��!���Z�c�*�5�x   x   ������m��2%�n�8�0�c�e~��ث�+�ϻ.������($��d7��'H��4U��]�=W`��]��4U��'H��d7��'$����M���C�ϻ7ث��~��:�c���8�Z%�x   x   �-���,��É�y%�&�5���Z�L����ʝ�����ڻ���BX�R���'��#0��4�ݗ4��#0�*�'�D��#X�����ڻ^���ʝ�4���b�Z���5��%����x   x   �l��*��R)���E��l���QŬ��ϻ�j����o;%� n9�/*K�sY���a���d���a�fY�)*K�n9�p;%�u��j���ϻ~Ŭ�P����l���E��Q)�x*�x   x   $'����,�U�A�qV]�����z��N���,�ʻ�
黒��&��'��N,&�=�*��*�&,&�B��.������
�1�ʻ����z�����RV]���A�9�,����&�x   x   �I)���,�PH3���<���J���]�vw�T(��N��ﰻ��Ļ�ֻ�����s��ֻ��Ļﰻ6N��Y(���w�@�]�
�J���<��G3���,��I)�#(�x   x   ,�E�H�A���<�T�8��A7���9�9�A�� O���`���u�p���S���OR��)���ℛ��Q��m���ȿ����u�e�`�< O�B�A�#�9��A7��8���<�ժA���E���G�!�G�x   x   �l�B]���J��97�!�%�u�����j�
����kO��"���'�j�)�B�'�n"��N�[��<�fj���������%��97���J�nA]���l���v��z���v�x   x   %������]���9������<���nD���en�Ikb�2?_�Y_�[_�B>_�fjb�Jgn�A���mC�� �����Y����9���]����O��晻N��������晻x   x   ᮬ��f��[�v�ϴA��������@|g�wQԹ-F=�Q~Y9��9��9�M:���9"��9�{Y9�!=��RԹ�}g����W���A���v�lf��ꮬ�C��8N˻�yϻ�M˻7C��x   x   vcϻ����/����N�TO��!���Թ�9�B:���:��:[�:�Y�:��: �:��B:m9�Թ� ��O���N���������cϻm뻗E��U��v���E��c�x   x   `H���ʻ�2���`�5������mS9�iC:ZA�:���:W�;~�;C�;-��:y@�:4C:r:9����������`�53����ʻeH���Q��e�:'��b*�+'��e��Q�x   x   �����軛ϰ��u�	s���m�;�Z9��:���:'�;ى!;�!;��;���:3�:)�Z9x�m�)r���u��ϰ���軞�� .)��.>�|DM��%U��%U��DM��.>�.)�x   x   �$%�P���tĻ��������a�pe�9�(�:��;i�!;��*;t�!;��;(�:�`�9��a�6 �4����tĻ(���$%���D�!�`��sv�(��Hz��5���sv��`���D�x   x   vU9�<��'kֻ������!�4�^�-��9N��:+�;!�!;��!;֑;Q��:���9&�^���!������jֻU���U9�� `������n��x����y���y��i����n������� `�x   x   JK�7���h1��u�'��\^���:��:~�;��;Z�;k��:�:0^^�M�'�1��p��I�-K���x��%��g!��%���"f��(���>f��#���;!��x%����x�x   x   ��X�	&�*a�/d��5�)��\^�}��9�0�:�
�:N
�:z1�:c��9o^^�@�)�d��>a� &���X������y�����ޝ˼�ټC�/��ټ��˼ ���y������x   x   _�a�R�*�����d��۝'�|�^��}�9�*�:�\�:.+�:{�9\�^�!�'�
e��	��!�*�l�a�q��0����Ǽ�V���5���g�G�����pV��ǼI���j��x   x   E�d��*�}d3��A�!�9�a�m0[94C:"4C:/[9��a���!��3��d��*�~�d�.���_ǲ�^�Ҽ���"���x�7�7��x�&�����b�ҼUǲ�?���x   x   �a��&�l�仑���#�X�m�r/7�B�9�:7���m��#�z�������&��a����(:���ؼ����1Z�s�����"����q�5Z������ؼ':�����x   x   ��X�����qֻߦ���u����Z�ӹ�ӹv���bu�Ʀ���qֻ�����X��!��fɲ�Y�ؼsf���i�Q���&)���.�Ó.��&)�G���i��f��l�ؼCɲ��!��x   x   �K�Ц��|Ļ��u�_�����ADg�������_�u��|Ļ���K�T������Ӽ�����j�N!�3.�͌6��k9���6�3.�[!��j�����Ӽ-���D���x   x   �]9����ذ�C�`��O�(�������O�]�`�ذ�g���]9�Y�x�=��ԼǼH��\�;��"4.�(K9��?��?�6K9�4.�1���\�V�𼳼Ǽ6��m�x�x   x   �-%����U;��b�N����j �3����N�`;����軻-%��+`�,��'
��c^�����))��6��?��
B��?��6��))����`^�=
��,���+`�x   x   g���ʻ�����A�������ùA�N��t�ʻ��0E��Ɓ��)��@�˼���}�����.�3o9�9?�-?�5o9��.�����}���K�˼�)���Ɓ�aE�x   x   �Y��Ò���v���9�_�%�.�9�	�v�&����Y���9)���`�yw��j�����ټk���n%��"�;�.�W�6��N9�d�6�6�.��"�w%�������ټl����w����`��9)�x   x   5sϻ�p����]�-:7�0:7�W�]�^p��4sϻ�\�=>�V�v����3r���%�{�j&����Q-)��8.��8.�E-)��r&�l��%�:r�����E�v�!=>��\�x   x   �������;�J��8�0�J�H������/,�s�;UM�Z'��΅��ò��'�����̀�&�j���#!�j��$�À�����%'�Ȳ��Ņ��Q'��jUM�s�,�x   x   ����HO]���<�	�<��N]�����)T��]��t'��8U�����놠��t���ټ��󼌠�Sb�Gq�Iq�_b����¬�	�ټ�t��������8U�5'�]��T��x   x   ��l��A��K3�5�A���l�3���Zb˻���s*�H:U�Y)��M�����v�˼�g�˘�&����u�����Ø�g�f�˼���Z��C)��I:U��s*���b˻"���x   x   l�E�y�,��,�V�E�~�v�˹��4�ϻ�	�# '�.ZM���v��|���0��h����ǼӼ��ؼ�ؼӼ��ǼT���0���|����v�?ZM��'��	��ϻ)�����v�x   x   �R)���OS)�?�G�� z�T���Ye˻�c��#x��D>��`��́��4������G���ײ�I���ֲ�K��������4���́���`��D>�Ax� d���e˻]���( z�V�G�x   x   �+��+�<'(�+�G�)�v������Z��/6��c�cC)��E�`;`�=y�1̆�&.���
���
��).��2̆�-y�B;`��E�eC)��c�6뻊Z������_�v���G�Z'(�x   x   �6���>��tY��т�����ɻl���\�v�7��XY��{�G7���������`E������mE���������K7���{��XY���7�\�����ɻ᧡��т��tY���>�x   x   ��>�0J���`�H���1���4��� ٻ�L�2���C1�n
J�$!a���t�<k��I'��8'��6k��Ϧt�!a�m
J��C1�"���L�Xٻ����ఘ������`�0J���>�x   x   hY�C�`�+n�����Ս��c��Uյ�^ѻ�𻎡��=(��.4��<���>��<��.4�5(�-�����ѻ;յ��c���Ս�����Dn�=�`��gY��V�x   x   qƂ�e�����������}҂��\��呻h}��mq��@mûˌֻ���F���a���X���I������،ֻ3mûeq��N}��呻�\��U҂�P�������ɤ��eƂ���������x   x   :������ʍ��̂���r�qe��_���a���j�!�x�vt��%ԋ�����uǒ�e���9ԋ�ht����x�A�j�ӷa��_�*qe�֭r��̂�Xʍ�ԡ��핡��k��t���k��x   x   S�Ȼ椵��Q���O��&de��,@���"���#`�����R���Dm�������zm������<���P`�h����"��,@��ce�P���Q��������Ȼ׻F�޻v�޻�׻x   x   ����� ٻ뻵�ё�ʌ_���"�-������(�|��Eu���Hv���8�/u�|v��0��g(�G����-���"�<�_��ё������ ٻ���	�g)����c)�=	�x   x   �F��9�D�л�b��"�a��r�����y�i����9��v:Jm�:��:��:�l�:2�v:��9��i�m���Gr���a��b��\�л�9��F�*�+��9�pA�!pA���9�-�+�x   x   m�7��q���P��f�j�m;�;�'�"��9:��:��:�_;p;�_;��:>��:u��9ݺ'�j;�0�j�5P���ﻝq�e�7�W,S�2�h�(�v�C�{�B�v�"�h�I,S�x   x   z:Y�J(1����Eû�x��������Fw:��:��%;\-:;<-:;Ѐ%;��:KGw:L��������x��Eû߉�b(1��:Y��~�c��@���������H���w��|~�x   x   q~{���I����`ֻLQ���f��������:�n;�3:;� G;�3:;�n;u��:���jf��^Q���`ֻ����I�j~{�-]���!���d��&�ļ�Pȼ6�ļ�d���!��=]��x   x   i$����`���'�;}�'����������@�:�/;�7:;8:;�/;
A�:�$��+���*���%}组�'���`�k$���J��SƼ%Oܼ�V켎��������V�BOܼIƼ�J��x   x   ������t�4�x��+͐�=���8�D�:Nu;��%;Iu;;E�:{8����=͐�x��44���t������b���{�q����*
��n�	���n��*
�X���	|༞b��x   x   ��vY����;����"��������K����:�9�:m9�:&��:������󟒻�����;�xY����2!мh���_ �-��(�c�-�k�-��(�$-�k �S���.!мx   x   1�����T�>������ΐ�x���p��rw:˩:|rw:-%��X����ΐ�����h�>����1���*ܼg��>����-�>�<�S~F�#�I�L~F�A�<���-�3��r���*ܼx   x   ���������;�l|�����Eg���ߨ��R�9�R�9ި�g������Y|����;�������Ow��
���#��:�};N�&\�cpc�gpc�"&\�y;N� �:���#�ױ
�Qw�x   x   13���[��K4�Ѓ绱T��������'�uvh���'������T�����{4��[��'3���x�/����(��>C�5�Z��m�A�x�D�|�>�x��m�6�Z��>C���(�=���x�x   x   t�����t�b(��hֻ��x�q8�Ɍ��&���B8�j�x��hֻM(�Њt�s���u.ܼ��
���(��F��;a�I�w����f`��g`�����K�w��;a��F���(�y�
�r.ܼx   x   *����a�d
�6Nû�j��k����k���j��Mûo
��a�3���I'м�����#��@C�D=a�V�{�9!��������������8!��P�{�D=a��@C���#����<'мx   x   �*����I����W��L�a���"�	�"���a�X������I��*��]j��%���ٵ���:�8�Z�Y�w�"���䐽�y���y���䐽"��X�w�=�Z���:�ʵ����uj��x   x   ��{��21����Ti��v�_�L@��_�Zi������21���{��S��v��D��-��AN��m�u�������z�� ͗��z������v���m��AN��-�O�}���S��x   x   �HY��{���л�֑��`e�`e��֑���л�{��HY��f���Ƽ�����4�H�<�A.\��x��c�������{���{�������c���x�C.\�G�<��4�Н���Ƽ�f��x   x   7�7��B�kƵ�dS��k�r�lS��PƵ��B� �7�.~�x-��K]ܼ3
��$(��F�Mzc���|��d��g���\琽b����d����|�Nzc��F��$(��2
�]]ܼs-��.~�x   x   S�[ٻ6Z��*΂�\΂�AZ��=ٻS��=S������r���g�Sx��-�l�I��{c�R�x� ���%���%�� ��V�x��{c�f�I��-�Wx��g��r�������=S�x   x   �������/э�ݞ���Ѝ�;���������+�i�y���I�ļ�������D�-�ƊF��2\��#m���w�9�{���w��#m��2\�ΊF�C�-��������D�ļ����i���+�x   x   	ɻì��l�������Ѭ��ɻ�	�x:�	w������bȼM���_z�w((�}�<��HN�
�Z��Ga��Ga��Z��HN�y�<�t((�fz�Z����bȼ�����w��:��	�x   x   Ԥ��J���6n�I�������j2׻9�݄A���{�Ꮯ�G�ļ�l��6
�+:�K�-���:�iKC��'F�lKC���:�P�-�*:��6
��l�1�ļ������{�߄A�9�R2׻x   x   zт���`�W�`��т�a}����޻��t�A�w����Px��xeܼ����S�m����#�	�(��(���#�i��S�����meܼhx������w�r�A���޻V}��x   x   �vY�Q7J��vY�>������\�޻Z;��:�x	i�Z���?5��Ƽ����������
�ܺ��
����������Ƽ<5��A����	i�	:�O;�L�޻���@���x   x   �>��>�;W�R����~���6׻	���+��GS�.<~��o���_���x��8м}Aܼ��⼏��uAܼ�7м�x���_���o��=<~�HS���+��	��6׻�~��c���\W�x   x   �5f�".s������'�ۻf���U0��	[�T����p���乼GӼi��'q��tb�U�jb�-q��h��GӼ�乼�p��S����	[��U0������ۻ����B��/.s�x   x   �&s�O#���g��]���GbѻL������&;��>_��҂�_������2��rC¼ȼ"ȼ�C¼�2��u��\���҂��>_�';�V�� ����aѻ߯���g���"��'s�x   x   �	���b���e��8���}�Ļ?��z(����1���K���e�J}���� 4���U���3�����@J}���e�n�K��1�+��N(�����Ļ;���9e���b���	������x   x   f����������ﷱ�aj���FĻ�*ֻ����@����[A$���1��<�H�A�]�A��<���1�)A$�����@�����*ֻFGĻGj������-���᢭�R���T񭻐�x   x   Q�ۻxLѻ��Ļ�a��{��層zԨ��I���x���Żk�ӻ� ��G�*.뻇G�r ໫�ӻ5�Ż�x���I��^Ԩ���z���a����Ļ^Lѻ��ۻ����I廼��x   x   �������C�ứ4Ļ�娻@��!※�k�d�`���]���_�(c�ue�due�;(c���_���]�_�`�Φk�!※����娻�4Ļ0��u���(��/��˹�ѹ���x   x   =0���	�uֻ{����؀��?�;m��ͺ�(���q��2M�ÝA�x3M���q��(��;�ͺqm�B�?��؀�����zֻ��P��==0�hFA��/L�u�O��/L��FA�x   x   ��Z��
;����@��-��n�k��[����0����:�J�:�d�: f�:bK�:)�:�4�����[��k��,��(�����
;�<�Z���u�Ą�!뉼뉼�Ä���u�x   x   '|���_�o�1��(�oS���T`���ͺ�R���׌:���:@�;�D%;k�;���:%،:'W����ͺ�S`�sS���(�K�1�n_�)|����X��\A�������A���X��f�x   x   Z��Y����K�r��M�Ż��]�Ι��<:���:'�3;	P;N	P;��3;���:�;:͙��]���ŻJ���K�e���Z���ɹ��м/"�4��	��"��м�ɹ�x   x   �ʹ�������e�S!$���ӻ�_���p����:�;�P;��a;�P;\�;ݒ�:P�p��_���ӻ]!$�§e������ʹ�ܼ�`���	���n]�"���	��`��!ܼx   x   �*Ӽ�駼 }��1���߻a�b�a>L��:"_%;�P;�P;5_%;��:V=L���b���߻��1�- }��駼�*ӼD���ƭ�f0#�/�<V5�5V5�
/�q0#����-���x   x   ��鼒�������;��/e�/�@����:��;C�3;��;���:?�@��e����;����~�����Ɍ��('�H�<�3�M�o�X���\�\�X�/�M�L�<��('�Ȍ�x   x   �R��
)¼���haA����e��5L�E��:�:c�:���:�3L�re���caA����)¼�R�����A)9��eT�2k�F�{�������U�{��1k��eT�<)9����x   x   AS�ȼ@���bA�5���b���p��u:��:Fu:�p�9�b�)軎bA�&@��%ȼ?S���$��@G�d	h�Cw��Q̍�G������6��T̍�Iw��Y	h��@G���$�x   x   �F�kȼ�����;��߻V�_�2���i�������F���^�_�R�߻t�;����dȼ�F���)��=P�*v�{�����������������������}���&*v��=P���)�x   x   �T��,¼T���&�1���ӻׄ]�Ƌͺ�~���ͺ_�]�H�ӻ�1�i����,¼�T���)�KUS���}�<񒽡�������d��<n���d���������7񒽫�}�bUS���)�x   x   �X����C)}�\'$�q�ŻfR`�2J��I��Q`���Ż�'$�/)}����X����$�9@P�4�}��%������ ɺ�,ǽ/ͽ%ͽ$ǽɺ������%��(�}�2@P���$�x   x   
����`�e����X���{k�]�?��|k��X����C�e����鼷��aEG��.v�󒽯���:����,ͽ�׽9xڽ�׽�,ͽ,�������󒽣.v�gEG����x   x   5Ӽ�����K�2/��0��'Ӏ��Ҁ��0��J/���K����5ӼԒ�09��h�􊌽����T˺�>.ͽ�\ڽ>� >Ὗ\ڽE.ͽ[˺����������h��/9�ے�x   x   �չ��Ƃ�)�1�w���¨�r����¨�f���1��Ƃ��չ������0'��nT�|��l!��z����ǽ�׽t?ὸ��t?Ὅ׽�ǽx���j!��|���nT��0'�����x   x   %e��(,_����_ֻ�䨻�䨻rֻ���),_�&e��a"ܼ�����<��=k�|ҍ�0����j��_�ͽa|ڽ�@��@�g|ڽV�ͽ�j��:���ҍ��=k���<����e"ܼx   x   ����5;�Z��;Ļ�w��R;ĻL�@;������׹��r��F;#���M�V�{����I"��yu����ͽh׽�`ڽZ׽��ͽ�u��F"�����Z�{���M�F;#��r���׹�x   x   j�Z������ỳe���e�������O�Z�� ��м�&	��%/�4�X�(������v#��/m���ǽ�3ͽ�3ͽ�ǽ&m��n#������(��/�X��%/��&	��м� ��x   x   �M0�������Ļ������Ļ�����M0�@ v�Dh��K6�a���d5�,�\�)���������A����Ѻ������Ѻ�A����������)���\��d5�g��M6�Sh��' v�x   x   ��]ѻ%���M���e]ѻ���ZA��ф�fS��ö�
k�f5�6�X���{�i֍��&��X�����������T����&��i֍���{�D�X�"f5� k����dS���ф��ZA�x   x   H�ۻ$���k��篭�(�ۻ����FL�����i���c�輞���)/���M��Ek�������������.��������������Ek���M��)/������{��������FL����x   x   �����k���k��п����⻁���P�����_V��g;༡*	�LA#���<�ryT�qh��=v���}���}��=v�~h�yT���<�@A#��*	�|;�3V������&P�j�����x   x   ��\(���������e廈��JL��Ԅ��m��/м�}��*���:'��;9�{SG�&PP��fS�5PP�|SG��;9��:'�8���}��м�m��Մ��IL�k���e廯��x   x   �1s��1s���������⻪���`A�
v�����Ṽ0ܼ&��d��5���%�?�)�@�)��%�4��m��*���/ܼ�Ṽ���	v��`A������⻸�����x   x   ����4��/����S��j���?� du��&��ׯ����������ws)��6�j3?�e"B�W3?��6�ys)���� ����ɯ���&��du���?��j��S�߹���4��x   x   �/���n���M����续���/�H�X�Qk��O����N�ؼA}�!�_�y�����_��C}�N�ؼ��	O��_k����X���/���^��QM��n���/��x   x   l����E���һL%�`���A��/9�*`Z�(��V������h���3�Ƽ��ϼeӼa�ϼ;�Ƽ�������P���&��M`Z�]/9�QA����8%뻫һBF����������x   x   �<���&�^�� ���c
��;�FG,��B���Z��+r��`��7 ��Z��c��P ��v`��\+r�ȣZ�#�B�4G,��;�fc
�&���1��%��绠<滕�����x   x   �X�N����������c�ʥ���Q�=u
��w�0� �Z)*���0���2���0�5)*�b� ��w�u
��Q������c��������?��c�cX�ڢ��&����x   x   ��?���/�,/�3V
��V��Wֻ`m»�Ӷ��|��PK������V��6�������V�������J���|��AԶ�qm»Xֻ�V�kV
� /�k�/���?�'�K���Q���Q��K�x   x   
Au��X��9��'����!`»�ʗ���n�J�?�� ��2�����]��;���2� �"�?��n��ʗ��_»����'�=9�`�X�Au�V����?��Ï��?��q���x   x   v��9W���=Z��+,��=����rxn����+�l�,#c�J� :o=F:X>F:�� :>!c���l�#��vxn�ߺ���=��+,�/>Z�=W��R��ow���ҹ����������ҹ�pw��x   x   K���x6�����}B��Z
��W����?���l���%:pL�:{;?�&;A;�K�:��%:&�l��?�W���Z
��}B���u6��E���9�ؼs�����r= ����~���ؼx   x   =�㼺ӻ�����1{Z��W����m����Y� m�:$);;w�`;o�`;�);;�m�:"�Y�������KX�4{Z������ӻ�E�㼘��A�n����%���%�[��A����x   x   n����ؼ�����q�d� ��r�����3k:�);L�`;N2x;9�`;);ol:����r��E� ��q�������ؼr���	�2�3���D���O��pS��O���D�1�3��	�x   x   /���Y�P����G���*����'0��#G:A�&;��`;�`;��&;�$G::0�����*��G��j����Y�(���B7�V�S��sk�)�|��ڂ��ڂ�+�|��sk�O�S��B7�x   x   �])�X�ŤƼ�押�Y0��h��=����2G:�4;�@;;b4;�2G:���Sh��dY0��押ǤƼK��])�3�N��*r��ш��-������˟�����-���ш��*r�.�N�x   x   ��6��K���ϼ��4�2��h���-���:-��:���:��:�-��h����2��񎼾�ϼ�K���6��b�����pT��h窽�ض�������ض�\窽nT�������b�x   x   @?������Ҽ�򎼑[0��������U�Cu&:;:U����&��>[0��򎼕�Ҽ���<?�tp����O먽�ｽeν��ؽܽ��ؽ
eν�ｽM먽���~p�x   x    B����I�ϼU銼�*��t��/��+l��+l�����t��;*�c銼Y�ϼ���B�wvw�H����e����̽H�὎#�$��'���#�F����̽�e��E���ovw�x   x   �?��N���Ƽ�K��� ����۠?�����?���Å ��K����Ƽ�N��?�xw�x���฽�9ֽ+��w���]���
��]�t��*���9ֽ�฽|���ww�x   x   J�6�n
�)���Cr��\�W��bn��an��V��!]�zr�"���r
�P�6��p�.����ḽ�wٽ`=�����g��'k�#k�e�����`=���wٽ�ḽ4���p�x   x   d)�d�����t�Z�3_
�����?�����_
�X�Z�����d�d)�b����Ai���<ֽ�>���
�5�#L�Ϲ�)L�5��
��>���<ֽ>i�����b�x   x   ���R�ؼꉓ���B��@��Y»�Y»�@�ՇB�����[�ؼ���7�N���������̽���^���5�b��x�#�v�#�_���5�b�������̽�𨽧���-�N�x   x   ����߻�H���4,�����YNֻ�����4,�1���߻�����L7��6r�2[������W�ή���N�|�#��&�}�#�N�����U������3[���6r��L7�x   x   ��B�� MZ��.��V�W�.�MZ�%B����k�{�S�tو��諾nν�,�4b��n�ȼ���#���#�Ǽ��n�1b��,�nν�諾qو���S�i�x   x   £���a��"9��[
������[
�"9��a��ʣ��	����3���k�87��U㶽��ؽ ��˒
��o�P�d��P��o�Ғ
� ����ؽX㶽E7����k�~�3���x   x   h����X��9�=���5����9�	�X�[����ؼ�M�~�D�2�|�����&����ܽ�!��d�����9��9�����c��!����ܽ'�����&�|���D��M���ؼx   x   PYu�Q�/����������/�xYu�������A��8�O��傽�ן�](����ؽ�1�%�����

����'��1��ؽW(���ן��傽A�O�:������x   x   ��?����'뻡'�����?����湼+���U�%���S��悽!��0綽�sν���E��]J��`J��?������sν-綽!���悽��S�I�%�9����湼.��x   x   th�m��qһ��ih�:�K��P��<����K ���%�m�O���|��;������������̽;Hֽ�ٽBHֽ��̽���������;����|�\�O���%��K �#����P��B�K�x   x   �S��R��rS��4T�T��J R�SՏ�����C���ض�X�D�]�k�c߈��b�����ft��xmct������b��Y߈�V�k�m�D����������Տ�. R�Y��x   x   �����u��񻷻�滭:��R��R��빼�~S���3�l�S��Dr�Y�������ʗ�N���ʗ����T����Dr�{�S���3�iS��=빼�R��R��:���x   x   R7���7�������i����K�
��c�����ؼ9���aY7�x�N�) b��0p��w��w��0p�4 b�t�N�\Y7��@��ɷؼ_���
��
�K�����滳���x   x   P��o�Ȼ��b��n�E����������nԼɯ�HM��;�W��Bo�p1���T��Zs���T��q1���Bo�#W��;�FM�����nԼ��������X�E�;�����Ȼx   x   ��Ȼ�ٻp=���
��S>�vn�气��7����ݼA���f���+�40<�_ H��kN��kN�` H�"0<���+��f�8����ݼ�7�������un��S>��=��x�ٻ��Ȼx   x   k���2��U5
�L���5�{�V����n
���1��v�ϼ�켪����Y�����J��'������켅�ϼ�1��m
��<��Z�V���5�.�p5
�`3��4��A�x   x   p�����Qx��)#�D.���>���U�4jr�Sԉ� ���$���۶��/�Ƽ�̼�̼.�ƼŶ�����1���Rԉ�jr��U�A�>� D.��)#�=x�Y�����&�;�x   x   Y�E�j>>�N�5��;.���)��h)��.��/9���G�D�X���i���w�O���N��e�����w���i�t�X�[�G��/9��.��h)���)��;.�m�5��>>�5�E��'K��M��'K�x   x   v|��fVn��V�$�>��_)��\���k��S�����f�$��4�����+��If�g��C����� ���\��_)�v�>�!�V�Vn��|���!���4���4���!��x   x   Ll��8���f��:�U�\�.�����6�?���\���I��ʁ}�~�q���m�Ѕq�*�}��I��']���>��q6����l�.�5�U�
��\���Tl��;b��{���Wüw��=b��x   x   \OԼ�����TDr�9����K.��7Yo�ڱ
��
���>��6��=r�k@��
���
��Xo�g.��
��89�3Dr��򗼎��SOԼV�����72�.2�����h�x   x   t����ݼ�������R�G�վ�5=��}�
��ȸL�:��
;�7;��
;�J�:�ȸ8�
��=�������G����������ݼg�����$��.��=1��.��$���x   x   W6������ϼl����X����|�����<x�:@m8;�*i;*i;m8;�y�:����b�������X�l���ϼ��U6�]�8���N�cR^���f���f�WR^�ÕN�W�8�x   x   ��;��O��뼁���6�i�=A�}��$����
;i:i;�&�;O:i;4�
;n!���}�DA�-�i���������O���;���]��{�l���bd��}��gd��p����{��]�x   x   +�V���+��������P�w����q�ֈ��g;�Ci;MDi;�h;��(q�6��j�w��������ͮ+�2�V�M�Gؔ�>���d�����������a���3���Oؔ�W�x   x   �#o��<�	����Ƽ����Ԛ��bm�;���D�
;}�8;��
;a���am��������ڙƼ
���<��#o�����;̪�P����MҽScݽi2�Qcݽ�MҽT���-̪�����x   x   �!��bH�t��q̼�2����q�ڹ�����:)��:����#q�,���2���q̼t�aH��!���ß����ٽ�?�� ��[��[��� ��?��ٽ$���ß�x   x   9E��'QN�)���r̼4���[���}��u��Y¸Jw���}�o�������r̼,��/QN�6E���婽 ,ͽ ���x������j����y������+ͽ�婽x   x   Jd���RN��u�Q�Ƽ:�w�C����r
�0r
�X���B�w�w�p�Ƽ�u��RN�Jd���5��g�ֽC���/��uT��)�\/�\/��)�xT�+��:���q�ֽ�5��x   x   �F��=	H����$����i����G4���(o�4����ՙi�������;	H��F���6���ڽ���>�v)��6�"�?�M�B�#�?�	�6�w)�>�����ڽ�6��x   x   �$���<�u��O��� �X�7�� ��V ����.�X�Y���x���<��$���詽�ֽ͹�H��3.��??�	dK���Q���Q�dK��??�3.�F��͹�)�ֽ�詽x   x   -o�V�+�E켂s����G�����"������G��s��7�Z�+��,o��ȟ�11ͽ����?�4.��B�znQ�[��n^�[�{nQ��B�4.��?����#1ͽ�ȟ�x   x   �V�<X�
�ϼ�É��9����Y���9��É��ϼ<X��V�4���Z�����Ȝ��)�>B?��oQ�W^�	e�	e�W^��oQ�>B?��)�Ɯ����d��)���x   x   e�;����p ��aQr�ۘ.��V��.�VQr�b �����i�;������Ԫ��ڽ#�eY���6��gK��![�z
e��lh�z
e��![��gK���6�eY�#��ڽ�Ԫ�����x   x   B�a�ݼ}���;�U��`)��`)��U�����l�ݼB�ޜ]��ᔽT����K�ء�k�)��?�ƸQ�s^��e��e�s^�ȸQ��?�k�)�١��K�Q����ᔽڜ]�x   x   ����*��ǝ���>�)���>�ǝ��*�����[�8���{�Ԛ��6[ҽ��1���c/���B��Q�o$[�<[^�x$[��Q���B��c/�0����B[ҽΚ����{�e�8�x   x   dcԼ����k�V��A.�vA.���V�����^cԼ���N��ˉ�����rݽ1d��s��d/��?��kK�uQ��tQ��kK���?��d/��s�1d��rݽ�����ˉ���N���x   x   �}���ln���5��-#���5�hln��}���#�q�$��g^�pq��I���C�e�D����)�I7�^H?�OB�`H?�L7���)�A��e��C�I��pq���g^�l�$��#�x   x   ��8P>�M��X��uP>�Њ��w��z���.�G�f��������uݽ��ͥ��^�B&)�<.�
<.�A&)��^�ͥ����uݽ������?�f��.����!w��x   x   ��E���;
�����E��2��+��B�5R1���f��s��ߵ��=aҽ5T�(����H�g��	H�����(�6T�?aҽ޵���s����f�=R1�B����2��x   x   ����D���E��ޒ��AK�=G��2qüC�k.��l^��ω�ؠ�����{ڽ������������������tڽ���ݠ���ω��l^�e.�C�aqü8G���AK�x   x   d��)�ٻt���$M�(H�����3��r�$�ۯN�X�{�r锽�ު��*���?ͽ��ֽ�#ڽ��ֽ�?ͽ�*���ު�t锽D�{�ԯN�u�$�@�����H��$M��x   x   �Ȼ`�ȻE-���BK�$5��<|���,�|$�H 9�K�]�a���ȑ��՟�{����F���F������՟��ȑ�Z��P�]�X 9��$��,�H|��)5��!CK����,�x   x   u�ﻪ* �{��)E�����櫼�9�K�)�2�SbY�����'���펤�1ⱽ�k��^\���k��1ⱽ펤�0�������EbY��2�K��9༇櫼y���(E�җ��* �x   x   & ����� #��G��z�믞��Ǽ�������3��Q�z:l�7���6쉽�M��}M��1쉽8���z:l�uQ��3�������Ǽ篞�(�z�!�G�� #�{��:& �x   x   ȋ���"�1�3�LM�2�p�ʮ�������μ��������y"�S]4�r�B�L�K���N�T�K�{�B�N]4��y"�������ؙμ{���ή��C�p��KM�;�3��"�������x   x   �E�W�G��BM���W��h�j����A���良�����ּ�@�z*��	������	�v*��@���ּ�����良�A��x����h���W��BM�4�G��E�*D� *D�x   x   �����z�G�p���h�J�d�z�f��!p�a]��{q��M헼���C������^������B�����Y헼sq��^]���!p�f�f�G�d���h�N�p�޾z����rH��ds��fH��x   x   )Ϋ���������p���-�f��R�[�D��,?���?��D��,J��O���R�j�R��O��,J��D���?��,?�U�D��R��f���������b���!Ϋ�*����Ẽ�Ẽ%���x   x   �༣�Ǽ�i��/���p��D�i"����U���׻��ʻ�Ļ�»�ĻB�ʻ"�׻�U����!i"���D��p�/���i����Ǽ��Y��N# ��Q�X# �?��x   x   �5�ʶ���yμ�ե��J���?����wջ��\w�k����˺=������˺v��]\w��ջ�����?��J��֥��yμĶ���5�����{+�_�1�Q�1��{+����x   x   ��2�G������;����X��V}?��+6w������":H2�:��;�3�:��":P���6w��+�M}?��X��(�������X����2�WtK�V_�^�k���o�^�k�J_�VtK�x   x   �BY�H�3�j��ǻּ�ϗ���C�%�׻���;d#:�);)�g;��g;�);!g#:���B�׻��C��ϗ���ּ���B�3��BY��
|�'���@S���蜽�蜽BS��$����
|�x   x   vv����P��^"���H���-�I���ʻ�˺���:Բg;���;��g;R��:�˺�ʻ+�I�L������^"���P�yv��)������G��6�ƽ�8ʽ*�ƽ�G�������x   x   <����l�n@4�6����-~O�,3Ļ�B���;�g;��g;z;ZC��h3ĻT~O����0�s@4��l�F����창\̽���C��������C�s��h̽�창x   x   �y������<}B���	�`ܴ��R��H»e8����:�-);��:z8��zH»�R�Eܴ���	�7}B� ����y���?Ƚe}��P� �����3����#��P�V}��?Ƚx   x   ṟ��ى�էK�����9����R��1Ļ��ʺU�#:m�#:_�ʺ�1ĻйR��9�����ߧK��ى�q̱���۽W��W��
H%��0��s6��s6��0�H%�Y��W����۽x   x   �U��I;���N����O޴�I�O�T�ʻ<{�7)��m|�F�ʻJ�O�8޴�����N�E;���U��t�����"�#���7�"G���P��0T���P�"G���7�(�#����k��x   x   �G��/<��x�K�n�	��"����I�}�׻
w��	w�O�׻��I��"��u�	�z�K�2<���G��>#񽞌��-���E��Y��g�z�n�v�n�
�g��Y���E�
�-����B#�x   x   aX��S܉�7�B�����*�C�q �߶��V �]�C�����)�B�X܉�XX���$�6���03��N���f�y��M���H���M��y���f���N��03�.���$�x   x   ѱ�,���3G4�)�՗��~?����'���~?�՗�/�=G4�.���ѱ����{���13���Q��hm�{��������!���!������v����hm���Q��13�}�����x   x   ���v"l��f"�6�ּ�]��2?��\"�?�	^��>�ּ�f"�x"l������۽R��M�-��N�#jm�ރ������P���z���P������$ރ�jm���N�P�-�Q����۽x   x   ږ��� Q��������N��V�D�E�D��N���������� Q�ۖ���HȽS��B�#���E��f� ������_l��M˚�P˚�al��~��� ���f���E�>�#�Z���HȽx   x   �~��y�3�0���sߥ�^p��R�kp�oߥ�)���u�3��~������c����_�7���Y��y�����GR��5̚���5̚�HR�������y���Y�c�7���]������x   x   #SY�����μ�6����f���f��6��ڈμ��#SY�١��v̽eX�WP%��G�|�g��Q��K%��F}��"͚�͚�C}��N%���Q��t�g��G�[P%�gX�}̽ԡ��x   x   �2�G���w�������d�����w��1����2��|�W(�����J%��0���P���n�tM��,&��
T��o��T��,&��nM����n�	�P�ݚ0�H%����P(���|�x   x   �C�7�Ǽ����N�h�0�h�����N�Ǽ�C���K�ֽ��hW���U�'���~6�X<T�&�n�KS����������������OS��,�n�O<T��~6�*���U�pW��׽����K�x   x   �0�����s�p�U�W�i�p�ܩ���0༬��L_��a��J�ƽ�����?�4�6���P��g�Jy���ヾ��Jy��g���P�6�6��?�����B�ƽ�a��E_����x   x   �᫼�z�?OM�YOM�[�z��᫼��󼻏+�o�k������Lʽ����L��v�0�G�ƔY�ʫf��tm��tm�̫f�ĔY�G�y�0�J�������Lʽ����|�k���+����x   x   ���϶G��3�r�G��������3 �E�1�Q�o�*���.�ƽ[�\)�V%�ð7���E���N��Q���N���E�ΰ7�
V%�X)�[�2�ƽ%���F�o�=�1��3 �#���x   x   �)E�#�#��)E��Y�����Cc���1���k�je��]�����
^�@��>�#���-��=3��=3���-�5�#�9��^����]��de���k���1�Nc������Y��x   x   e����� ��BD�ǅ��$���Y5 ���+��#_�%Ì�0���(̽ܖ꽧��%����x�����'�������(̽0��)Ì�$_���+�N5 ����̅��BD�x   x   - �0- �����AD��Z��?�����󼪯���K�$-|���������WȽ"�۽����:��:���� �۽�WȽ�������3-|���K�������M����Z���AD�S��x   x   H����!��1C�w�|��
����߼P��*=�ISm�Bؐ�:���ݖŽ�iܽXU�\�������b���XU�jܽ�Ž4���7ؐ�LSm��*=�S���߼�
��i�|�2C���!�x   x   ��!���0���O�:��5V����μ�/���#�c�H�.-p��ߋ�zM���׭����������������׭�mM���ߋ�F-p�|�H���#�t/���μ<V��8:����O���0���!�x   x   Y"C�k�O��Mf�X��_k��	���q��	��+#�o�>�c�Y��;r�3ʂ�����'�����*ʂ��;r���Y�w�>��+#��	�r���Tk���W���Mf���O��"C�
?�x   x   b~|�:/���Q��b؋�旼tP��{���}9ݼ����`��!��/��#:���?���?��#:��/��!��`�����9ݼt���FP���嗼�؋��Q��9/��b~|��{�{�x   x   T���gC���]���ޗ�qJ���阼�m��ɤ���{���μm߼�G����q��������G�i߼�μ|��Ȥ��`m���阼�J���ޗ�~]���C��F���L���w��M��x   x   ��߼��μX����@���ᘼC������~���ك����ꕌ�<Ր�oH���H��KՐ�Օ��"����ك��}�����p���wᘼ�@��r�����μq�߼@;�r��T��/;�x   x   >����;Q㼞m���\������_�+�?�dL*��P�4F�2���.�&F��P�L*���?�P_�����\���m��PQ���@��9����'��*���'�(��x   x   �=�$�#�q��fݼ����Jn��b~?�-	�»U���Z�P��w0�*w0��P�t���5»^-	�N~?�n��񋬼�ݼq���#��=�asR�? b�F1j�71j�A b�gsR�x   x   �/m��H�#�����g[��.Ã��0*�X����+�����lbt:�`�:�^t:E���)+������0*�<Ã��[�������#��H��/m� ㆽ������۞������#ㆽx   x   Ð��p��>�zG���ͼ¢���*�:s��Ԇ���#;	JZ;4JZ;�$;r����s��+�΢����ͼ_G��>��p�Ð��ǧ��-���7ɽ,�н>�н�7ɽ�-���ǧ�x   x   ����ʋ�ʻY��� ��޼Mu�����gP�Aeu:�dZ;�;|dZ;`au:/gP���Lu���޼�� �ۻY��ʋ����CXʽ���5����L�����L�=������7Xʽx   x   :|ŽW6��Sr�j/����`��I�/���:�tZ;�tZ;P�:��/�n������
�j/�Or�N6��B|Ž�|�-8�j@��"�(�'�(�'��"�j@�/8��|�x   x   �Mܽr�������:�p{��$������/�O�u:DV;�u:9�/���$��m{���:�����v����Mܽ���Ԋ��d0���?�I�I�8M�O�I���?��d0�֊����x   x   _8� ���.��?������$������RP����	���RP�����$��������?�6%���[8�����A.�z&G�5�[�Duj��r��r�Auj�=�[�y&G��A.����x   x   ����f澽��ף?��}��w�����0a����*��a����u���!~��ޣ?����]澽�����K�%<��Y���s������1��{Z���1��������s�	�Y�!<��K�x   x   ����羽�:�%�=w��6'�����S���$'�Rw���:���羽*����0!��D�s,g�����ҏ�.ט�������,ט��ҏ����u,g��D��0!�x   x   ������U���`o/���޼Ƥ���)*�	��)*�Ǥ����޼ao/�X������ޭ���1!���G��n��舾�A������o��&����o������A���舾�n���G��1!�x   x   �>�$ŭ��r�w!�2�ͼ�ă��s?��s?�~ă��ͼ�!��r�ŭ��>��N�x�D�?n��㊾v���#���;���~���~���;����v����㊾Bn�s�D��N�x   x   OVܽq=����Y��N��b��	n���^��m���b���N���Y�u=��RVܽ����<��0g�9ꈾ`���xq��9J���V¾už�V¾:J��{q��^���4ꈾ�0g��<����x   x   �Ž�ҋ�y�>�6�������������񑬼�����>��ҋ�~�Ž���5H.���Y����eD����HK���ž"�ʾ"�ʾ�žHK����hD�������Y�9H.����x   x   ����p�:#��$ݼa��g���a���$ݼ?#��p�������ђ�0/G�|�s��֏�����>���X¾F�ʾ0U;F�ʾ�X¾�>������֏���s�,/G�Β����x   x   2ΐ���H����~x���㘼�㘼�x������H�4ΐ��fʽ�@��n0��[��惾�ܘ��t��,����žo�ʾo�ʾ�ž,����t���ܘ��惾 �[��n0��@��fʽx   x   �Dm���#�mc��H���J��I��Jc㼝�#��Dm��է�f��K���?�F�j�o8������8���F���>[¾ž>[¾F���4�������w8��B�j���?�K�h���է�x   x   � =�|(�:
���䗼�䗼C
���(�� =�3����>��m���8!"�F�I��+r�b�������v�� B���O���O���A���v������b���+r�M�I�>!"�q����>��2���x   x   Y ���μ$i���܋�i��s�μX �\�R�ғ�KɽY�6�'��+M�k-r�9:��vߘ����A���w��D�����tߘ�?:��n-r��+M�3�'�Y��Kɽғ�`�R�x   x   ��߼�S��^Z��mZ���S����߼n���b�!��E�н��h�'��I���j��郾�ۏ�J��������J���ۏ��郾��j��I�d�'���N�н#���b�c��x   x   x��t;���Yf�U;��z���Y�w�'��Nj���н�Z��$"�6�?���[��s��#��-��늾,񈾺#��"�s���[�1�?��$"��Z�۬н��Nj���'��Y�x   x   x�|���O� �O���|�6���L�*�WPj�o��Pɽ����P�7v0��8G�u�Y�p>g��$n��$n�t>g�i�Y��8G�>v0��P���� Pɽx��fPj�F�*���2��x   x   o5C��0�F5C��6{�<���Q���'��b��֓��E������G����'S.��<�*�D���G� �D��<�/S.�����G���彪E���֓��b���'�T�X����6{�x   x   ��!���!�x-?�p6{�a���]켾��%�R�W����ާ��rʽk��~��? �\�s@!�y@!�\�7 �~��n���rʽ�ާ�S���"�R�İ��]�\��C6{�Q-?�x   x   �;��%I�t�C����Լ�����<��8t��ܙ��Z��k�߽�� �{��F�'�"��8%�"�"�F����� �^�߽�Z���ܙ��8t���<����$�ԼG���Jt��%I�x   x   >I�Nj\�2.��i����ͼ�,�E�(���S�=M��pW��p���ν�	����n���n��"��	�ګνp���W��?M��b�S�2�(��,��ͼk���*.��'j\�-I�x   x   n�s�I(��LՐ�ZM��)�Ƽ���x�bl1�4)T���x�;X��/o���-���\��3/���\���-��5o��NX����x�)T�dl1�Bx�����ƼQM��RՐ�G(����s�e�n�x   x   4Ꞽm���lE��ǆ��������ټ���7��^�%�X�<�F*S��Yf�\pt���{���{�ept��Yf�=*S�H�<�e�%�P�����o�ټ��������gE��l���1Ꞽ����x   x   _�Լ��ͼ^�ƼT�������3{ż�zм5���a��z���/�Q���#�bV%��#�_���/�m��!b��9�Ἢzм<{ż����L���1�Ƽ��ͼj�Լ��ټK�ۼ�ټx   x   ���M�7��Coټ�pż]���Wh���G���-���G���v��t�¼+Ƽ-+ƼW�¼�v��)H��.���G��:h�������pż�nټ?��f����ר�������Ԩ�x   x   9�<�́(��b�޲��[eм�]��>ɓ�7����,h�B�Y�R�qO��=N��O�aR�.�Y�g,h�.����ɓ��]��2eм���c�(�-�<���L��UW�c�Z��UW���L�x   x   et�R�S�bP1���
|�p3������^�=��8�b#ջ3������������_#ջ9���=�����3���{�.��]P1�9�S�ft��Ƈ��Ǒ�h��h���Ǒ��Ƈ�x   x   �ř��8��eT�k�%��7�����l	h�)�r��L�ٺ+���bI�9����,�ٺr���(�?	h����#8��j�%�MT��8���ř�=Ʈ�}]���ʽ��ͽ�ʽ�]��>Ʈ�x   x   ?��?����x�3�<���b#���TY��Ի�^ٺ�λ:y1@;i2@;}ѻ:x_ٺ1�Ի�TY�u#��	���<���x�,?��?����ٽ3 �k��	H�H�j��( ���ٽx   x   �߽�T��A���S����L���Q�|Ϋ��n���R@;�Y�;�R@;����PΫ�'�Q��L�����S�A���T���߽.������"��+�x�.��+���"���,��x   x   q� �֍νV���1f�\���u¼��N������y�9�g@;�f@;nz�9)�����N��u¼P���1f�V��ˍνq� ����A�0��8D�XR��MY��MY�\R��8D�<�0����x   x   1���⽊���Ft���"�F�ż%�M�����7���L�:���P���j�M�F�ż��"��Ft������7��*&.�7*K��d�4x�[�����[��4x��d�A*K�(&.�x   x   Y3����>B��ټ{��6%�,�ż5�N������غ��غ.«��N��ż�6%�Ҽ{�=B����Z3�	�>�?�a��À��΍�1��웾웾5���΍��À�=�a��>�x   x   ��"�pO�����f�{�� #��w¼t�Q�*�Ի�C��A�Ի7�Q�x¼� #�f�{����jO����"�kK�;rs�I�������ǉ���u��f*���u��ȉ������H���7rs�iK�x   x   '%�Q���D��)Kt�Ϫ�cO��mPY�N��wPY��O�����Kt��D��Q�� '%�HQ�p�~����'��������þ1�ɾ4�ɾ��þ���*������n�~�HQ�x   x   ��"��������8f�Q��&��h�Ƈ=�Wh�i&��R��8f������񽻝"�oIQ��+���j���ٯ�þ��Ѿ��ھ-޾�ھ��Ѿþ�ٯ��j��,��sIQ�x   x   [7�w��\���S�
�����=���4������	���S�\��n��[7�CK���~�pk��eU��xȾ�nھ�羿�������nھ xȾgU��ok����~�BK�x   x   ɖ�#�νDH����<��A���3��9���x3���A����<�DH��.�ν˖��>�?xs�����ۯ�@yȾhgݾP\�Z�������Z��O\�bgݾ?yȾ�ۯ����Cxs��>�x   x   "� �_���x���%�V�Ἰ[���[��@���%���x�_��� ��-.���a��������gþ[qھ�]�f����� ��� �`����]�_qھfþ���������a��-.�x   x   h�߽#J��AT�٣�:kмԹ��-kмޣ�HT�J��i�߽���|4K�Jɀ�O���v�����Ѿ��U]��C� �)�C� �W]���羱�Ѿx���O���Iɀ�~4K����x   x   �M��=C��%^1�j���tż�sż����^1�9C���M������ 1���d��Ս�ǐ��A�þ*�ھ
�������� ��� �������,�ھB�þĐ���Ս���d�� 1����x   x   �ә�b�S�o�hzټ����vzټ�n�p�S��ә�\ڽ~+��FD��Cx�g ��(~��N�ɾ�޾b��.`������%`��d��޾N�ɾ)~��g ��|Cx��FD��+�fڽx   x   H,t�U�(�۪��������Ԫ�]�(�:,t�l׮����"�c R�d��y����3����ɾ��ھ��c�c����ھ��ɾ�3��{���d��h R���"���g׮�x   x   P�<�(�w�Ƽ}���n�Ƽ
(�K�<�և��q��\��Ŷ+��_Y��������]�����þ��Ѿ�wھoݾ�wھ��Ѿ��þd���~��������_Y���+�`���q��և�x   x   ����ͼ�P���P���ͼ�����L��ؑ��ʽkV���.�KaY��e��b#�����'���~þ��Ⱦ��Ⱦþ,������^#���e��MaY���.�mV�wʽ�ؑ���L�x   x   ��Լ����ܐ������Լ����qW�� ����ͽnW�?�+��$R�<Jx�2ڍ�a�������䯾C_���䯾����_��4ڍ�@Jx��$R�8�+�lW���ͽ� �� rW����x   x   �����2���2�������
ڼ���[��!��}ʽA��r�"��MD���d�Vπ��L��7u��7u��J���Xπ���d��MD�u�"�F��zʽ�!���[����
ڼx   x   �t�Xv\��t�����ۼ���tW�&ܑ��w����2�y	1��?K���a���s�-�~�:6��(�~���s���a��?K�|	1�2���w��#ܑ��tW�����ۼ��x   x   �)I��)I��n����ڼG��y�L�ۇ�T߮��ڽl�����t:.��?�2K�%\Q�-\Q�3K��?�x:.����n���ڽM߮�ۇ�w�L�I��ڼ����n�x   x   td�_�u�w����9ļu@��_2� m�L�� �½d����T#��6�޴D�@�M�2'Q�3�M��D��6��T#����\��5�½O���m��_2��@��9ļ]���U�u�x   x   ��u�+䆼����2�Ǽ���+%���S�������lsƽ7���V��A�Č��h��h�ˌ��A��V�E��|sƽ���������S�+%������Ǽ����H䆼��u�x   x   "������(����
ϼ�j����q98��5`�҅������-����ɽHڽ�~作��~�Aڽ��ɽ�-��v��؅���5`��98���ej���
ϼM���������{b��x   x   4#ļ��Ǽ� ϼD`ܼf��V�h���5���R�ۜp�P���M���,����������-��G��H����p���R��5�\���V�a��``ܼ� ϼ��Ǽ7#ļ��¼��¼x   x   I.�Y���T��F��={��u������[�a����-���<�mJI�N�Q�X�T�a�Q�yJI���<���-�h���[����v��g{�O���S��@���].�pR�)x�~R�x   x   �D2��%�Aw��I��h����%�ݼ�qܼ�bἪM꼘l��;��� �� �� ���l���M��b��qܼ�ݼ�缜h���I�9w��%��D2��@<���A���A��@<�x   x   n�l�^�S��8�������ݼ�y�����������\�����Ί����	]������������y����ݼ�����8�T�S�_�l�����3D��'���+D������x   x   ~�������H`���5�HG�5Xܼ���ݤz�?�Z%��4��O��}��#4��=%�?��z�����Xܼ9G���5�@`�����{��� G��A㷽"���/���<㷽G��x   x   ��½�򤽭o��8lR�����=Ἰ���0?���ٻI�W� ���nI�ŝ����W�n�ٻ:?�����>ἱ��DlR��o���򤽤�½�ݽ����b��� ��b������ݽx   x   i�Tƽk���rp�aq-�y꼠9�z�W��5�9�\;^;�;�9˝W����r�]q-��rp�[���Tƽo��v
����5"%� +�+�3"%����x
�x   x   ���@��?������/�<��7��_8��#����δ�څ;�8e;م;\д������8���7��5�<�����L��C�����D�&���<���M�N�X���\�V�X���M���<�J�&�x   x    ?#��C�ҧɽ����=#I������ꊼ݂�lwG�q�;.�;�vG�_�绾ꊼ����$#I�����ϧɽ�C��>#��B��_�ܝw�/g���㈾�㈾0g���w��_���B�x   x   � 6��-��ٽ����pQ��� ������}�0���ɑ�9*����}������ �"qQ�����ٽ�-�� 6��:\�*���ݏ���Oģ��i��Iģ����ݏ�*��{:\�x   x   y�D��x��]�U࠽rXT�&� ��ꊼ=����VW��WW������ꊼ� �kXT�G࠽y]何x��D�W:q�C���͡��ݱ�/I��8þ8þ4I���ݱ��͡�C��Z:q�x   x   (�M�U�+��QᠽksQ������7��,��[�ٻ����7�������sQ�JᠽG��U�"�M�j��&��Ml��twľM�Ӿ=�ݾ���3�ݾO�ӾzwľHl��%��m��x   x   Q�)V�t`�{���'I��;��9쏼�>���>�Z쏼�;���'I�z��o`�!V�Q�����B��������Ҿ)� ��������#��
)��Ҿ����=�������x   x   ��M��{���ٽ>���<��#�2���ևz�=����#��<�H����ٽ�{���M������M�����ǎ۾!�z�\��

�_��z��Ŏ۾����M������x   x   ��D�l2���ɽ5����w-�Aἁ���i���"A��w-�8�����ɽk2���D����.��������޾1���������͎�Ȏ�������7�����޾���,������x   x   6��I�t��?p���Yܼ|n��Yܼ��"p�~���I��6��Aq��!��ú�F�۾�����	�)b���M����(b��	�����L�۾ú��!���Aq�x   x   pG#�̻�$���xR��L���ݼ��ݼ�L��xR�*��»�lG#�AD\�MH���q���Ҿ5�h���b�����������b�k��0��Ҿ�q��JH��@D\�x   x   ����bƽZy��6�5�'��5�"��A�5�Zy���bƽ���:�B�v0��iԡ�S~ľ�/澡}�����������!����������}��/�Q~ľjԡ�y0��4�B�x   x   	��\ ��$`�n��cm��Im��{�� $`�` ����(�&� �_��叾汾��Ӿ]�� "���۝�������ޝ��� "�d����Ӿ汾�叾!�_�/�&�x   x   k�½լ��.8�Q��|�Q�.8�㬅�]�½;
���<��w����BS��p�ݾ���h
�ݒ�r�����k��ޒ�m
����f�ݾES������w���<�?
�x   x   g	����S�ڃ���*��σ���S�`	���,ݽ���5�M�)q��Hϣ��CþT��F!���#�U��Kf�Of�Y���#�@!��\�ྔCþDϣ�(q��:�M�����,ݽx   x   am�7%%�ag���gܼcg��F%%�]m�fZ��q�2%���X���u���Dþ!�ݾ��󾱀�Z����	�X��������!�ݾ�Dþ�u�����X��2%���\Z��x   x   �Z2�[����ϼ�ϼJ����Z2�����z������F&+�)�\��pѣ��V��#�Ӿ�6���ޮ��ڮ����6�$�Ӿ�V��qѣ��.�\�B&+����|�������x   x   �>�4�Ǽ����L�Ǽ�>��Y<�DV������S��'+��X��s������뱾ȅľ�Ҿ�۾��޾��۾�Ҿ��ľ�뱾����s�� �X��'+�a�����EV���Y<�x   x   �:ļk��Z���:ļ0e�e�A��������؃��16%��M���w��돾�ۡ��z���ͺ��$���$���ͺ��z���ۡ��돾��w�$�M�86%������������i�A�3e�x   x   "����놼.���7�¼�����A�X������������<�/�_��7���P���+�����1Z������+���P���7��9�_���<���������$X����A����,�¼x   x   K�u�C�u�Oq����¼)f�#]<�3����`���6ݽy#
��&���B��S\�STq�S%��*	��,	��U%��PTq��S\���B��&�|#
��6ݽ�`��/���]<�f���¼[q��x   x   I"���咼�㳼��-� �� Z�����~ҽ�{r����M/�֛I��`��Rr�O�}�����A�}��Rr��`�қI��M/����r�ҽ������ Z�D� ���4㳼�咼x   x   �ߒ�װ��+{���`�~��I�	���ä�g�˽,w��j�v"��W2���=�D�C�U�C���=��W2�v"�j�.w��R�˽�ä�	����I�~�\`�>{��+����ߒ�x   x   oԳ�r��TA׼q����c�X�7�w1b��3��IO��5�ý��-(���*�]��"��R���*�E(��֏��ýeO���3��b1b�Y�7��c�����vA׼�q��2Գ��ϯ�x   x   � ��J�������_*�"�&���@�'�`� V��%C���]��h嶽�D½cGȽ[GȽ�D½Y嶽}]��CC���U����`���@�-�&�d*����"����J� ��w뼊w�x   x   �� �k��U��"�g�PI�\Z"��S1���C��#X��~k�t�{�U��E焽g��v�{��~k��#X���C��S1�zZ"�\I��f��"��U�k�˨ �t�$���%���$�x   x   ��Y�,�I�9�7��&�A��"��	�j	�u���� �����#��#���� ���c��z	��	�u"�A��&�/�7�4�I���Y� *f���l���l�)*f�x   x    }����b�F�@��I"��	����@*Ѽ����8���1-���a��xU���a���-����������b*Ѽ��뼩	��I"�H�@�b���}�����U+������=+�����x   x   �����������9c`�~:1�w��qѼ����z��K��q0���#�p�#�=q0��K�%z�^���yѼ���q:1�c`��������ﴽ�&ӽ<�⽰�����9��ӽx   x   �M���˽�3���?����C����M�����y��H������K�E��>�K�:��AI���y�j��������C�@���3����˽�M�Kk�UB�U}�S �X}�RB�Lk�x   x   �w��P��ޯý)����W���\��5�K�K�z�b�Rb�:�d�:�b��𮻻�K��\��� ���W�)��ʯý�P���w��o*���=�'�K�	�R���R�*�K���=��o*�x   x   -5/�}T��k�3@���Qk�S��� ���90�5HK��ĩ:K�2;�ĩ:.HK��90�� ��i���Qk�'@���kགT�45/�J�M��vh��b}��X������X���b}��vh�T�M�x   x   ?�I��^"�� ���Ŷ�X{�����0��I�#����:���:��2�#��0������W{��Ŷ�� ���^"�5�I�6�o���������q��$ݧ�&ݧ��q���������6�o�x   x   "m`�W?2�'�G$½y�����"�^#����#��"K�,a�� K���#�U#����"�����P$½.�N?2� m`�3r���N��sF������-DȾ�s˾$DȾ���uF���N��0r��x   x   X6r��=�܊��&Ƚ�΄�e�"��0��f10��Ʈ�EǮ��10��0��h�"��΄��&Ƚъ��=�_6r�C(��ZN����ž�-پo���s�澿-پ��ž^N��A(��x   x   Hx}��C�<��!(Ƚ�����P ��H�K�(��K�" ��������(ȽK���C�Ix}��/��[��8c׾1{ﾞ������������7{�1c׾[���/��x   x   ����j�C�����'½�]{���bZ��G�y�h�y��Z��*���]{��'½���_�C������ߡ�^�þ����> �����H�^��]���H�����> ����V�þ�ߡ�x   x   f{}���=���w˶�!Yk������)韼������'Yk��˶�����=�u{}��ࡾ�_ƾ�'꾶��8��Ɔ��Z%�0�'��Z%�Æ�4������'��_ƾ�ࡾx   x   u<r�E2��
��?G��X�����Ѽ�Ѽ���$X�@G���
��
E2�x<r��2����þ�(꾊c����x�$�Z.�F;3�B;3�Z.��$�����c��(꾭�þ�2��x   x   �u`�f"��v��0����C�m��V��n����C��0���v�	f"��u`��,���_�����5��Ь�3#'��3��|:�m=��|:��3�,#'�Ӭ�:����㾍_���,��x   x   ��I��\��ý�G���A1��	��	��A1��G���ý�\���I�x���T��|i׾�A ����F�$��3���<� "B�"B���<��3�I�$�����A ��i׾�T��x��x   x   �@/�db��@��Mq`��N"�Y��N"�^q`��?��Zb���@/�� p��V����žm�ﾉ��C���\.��~:�1#B���D�0#B��~:��\.�A�����j�ﾵ�ž�V��� p�x   x   ����˽�(��X�@�<D�1D�]�@��(����˽��ܽM�#���P���7پ���M�v_%�6?3��=�D$B�F$B��=�3?3�u_%��M����7پP��$����M�x   x   d�����H#b���&�h���&�S#b�����c�(~*���h���r����澧��V��õ'�9@3��:���<��:�:@3�ǵ'�S��������{������h�)~*�x   x   �Ƚ�C����7��)��)���7�:���Ƚ��x��=��w}��}��`QȾ[��<��fa%��_.��3��3��_.�aa%�;�����`�WQȾ�}���w}��=��x�x   x   ҍ����I�b���
b���I�Ӎ��ӽLR�7�K��d���ꧾS�˾��H���P�����$��('�
�$�����P�D����T�˾�ꧾ�d��=�K�VR�ӽx   x   ��Y��{�ʒ�����{���Y����ͪ�R��D�R�����맾�SȾ����
��������������
�����SȾ�맾���<�R�A��٪⽶��x   x   O� �
c�bM׼4c�S� �If��A���꽍f ���R��f���������>پc��NG �����j����LG �[���>پ�������f����R��f ��꽹A��mIf�x   x   ��|���O������$��l������꽩����K��~}�U��W����žbt׾���R7�J7���ot׾��žW��U���~}���K�����������l���$�x   x   �泼�����泼c��`&�w�l� D��ɯ⽷V��=�ɒh�ڑ��*_��_���k��q�þ�nƾy�þ�k��_��/_��ߑ����h��=��V�د�	D����l�@&�N��x   x   �蒼�蒼⯼ǖ�ܝ$��Mf����$ӽ�~���*���M�Op������7��_?����a?���7������Ep���M��*��~��$ӽ��mMf�֝$���-⯼x   x   i螼Bǫ�^QӼ��"?��0��ܑ��>6佻��H�1���R��>r�=����B���藾|.���藾�B��:����>r���R�C�1����@6�鑮��0��?����PӼ8ǫ�x   x   %����u��M]�ٚ���8���p��ڛ��ƽ������H�,���C���V�:1d�4Ek�@Ek�81d���V���C�K�,������ ƽ�ڛ�o�p���8�ʚ�x]�Uv�����x   x   -?ӼNR⼛���C!���2�9m[����+���rȽ�P�X���� -#�9�*�,�-�1�*�)-#���R���P��rȽ�+������@m[���2�N!�����3R��>Ӽ�sμx   x   � ������!R��.�m�F���f�v��qS��G�����ʽћݽ�t�^��[��t�Ûݽ��ʽf���mS��\����f���F�+�.��Q����� �����x   x   ��>���8���2��.���/�� 6���B���U�#?m��;��hF��(9���Ɵ����Ɵ�"9��~F���;��?m���U���B�� 6���/�
�.�у2���8���>���C�NE��C�x   x   �����p�3Q[���F���5��u*��A%�H&�	�+�#(4��:=�U�D���H���H�H�D��:=�(4���+�]&��A%�hu*���5��F�3Q[���p��������������������x   x   [v�����m����f�@�B��7%����G����j��3漹�㼸�����´��㼣3��j�p�������7%�X�B���f�vm����ov�������eǽ�ʽ�eǽ���x   x   ��5�Ž-��S����U�&�q�����Ƽ^잼������k��^��^�~�k�����q잼��Ƽ����&���U�C��'��M�Ž�佑����4�U"�\"��4�����x   x   ����f���QȽ�8��$m���+��I��ݞ��L�6�K���<������5��L��ݞ��I�+��m��8���QȽ�f������$$��3�Ce=�P�@�He=��3��$$�x   x   m�1�*��*��g���#���4���䄼� ��4�(ǋ�q�����4�� ��ㄼ�漬4��#���g��*�"��i�1���L�}�c��t�G*}�7*}��t���c�y�L�x   x   ��R���,��|�d�ʽR+��|=�k~�o�k��������`ȷ:����Z���|�k�o~㼐=�e+��Y�ʽz|���,���R�'w��v���ᗾƟ��z��Ɵ��ᗾ�v��1w�x   x   1r�ĈC����uݽ���D��z�u�]��㕻�刹=䕻��]��z���D����uݽ��͈C�&r��㏾ˬ���ൾ',¾{�Ⱦ��Ⱦ&,¾�ൾʬ���㏾x   x   ����{�V��#��M뽵���j�H�����]�8���p!4������]���f�H�¨���M��#�t�V�����v/�����+oҾ���?����6���*oҾ���v/��x   x   2���d���*�w���F�H��z�Y{k���4	��{k��z�O�H���o���*��d�2���*��_о���;P��o	��������o	�8P����`о�*��x   x   ;ؗ��(k�r�-���򽠪����D�]~��ۄ��aL��ۄ�&~㼃�D��������x�-��(k�Aؗ��Ȼ��X߾Z4 �q��l��] �{�"��] ��l�q�W4 ��X߾�Ȼ�x   x   ���*k���*�
R뽔��=��漏О��О��(=����R���*�	*k�����I��{���x�x��f&��N0��u5��u5��N0��f&�x��x�s�辖I��x   x   ڗ�;d��#��|ݽ0���	4��D���Ƽ�D�~	4�0���|ݽ�#�7d� ڗ��J��]D�c;������/���<�j�D���G�l�D���<���/����e;�aD쾹J��x   x   �5��I�V������ʽ%)����+����������+�.)���ʽ���K�V��5��̻�0��,<�J� �%L4��5D�p�O��rU��rU�o�O��5D�'L4�E� �,<�0��̻�x   x   ������C�d���q��Q!m��&�����&�F!m�vq��d����C�����0��^߾{�y��#M4�=�F�*U��=^��Ya��=^�*U�8�F�&M4�}��{�^߾0��x   x   w+r���,��8�_B����U��6%��6%���U�eB���8콊�,�q+r�p6���о8 �w{���/��7D�=+U��@a�b�g�b�g��@a�?+U��7D���/�v{�
8 ��оs6��x   x   ]�R����c`Ƚ���B��q*��B�
��\`Ƚ���`�R��돾��S���u�:k&�ȉ<��O�@^���g���j���g�@^��O�ǉ<�:k&��u�U�����돾x   x   D�1�G{�������f���5���5���f����Q{��E�1��%w�����vzҾ5V��r��T0��D��wU��]a��g��g��]a��wU��D��T0��r�2V�rzҾ�����%w�x   x   ���ƽ8y����F���/���F�<y��ƽ����M�\���?����v	��d �}5�<�G��xU��B^�xDa��B^��xU�=�G�}5��d ��v	���A�\����M�x   x   �*佻қ�nd[�v�.�n�.�ed[��қ�~*�5$�Jd�=c:¾��������"�&~5�3�D���O�&0U�)0U���O�0�D�(~5���"�������_:¾:Jd�5$�x   x   ˊ����p���2�nW���2���p�Ҋ�����D�3��t�'ԟ�q�ȾS�򾧲��f ��W0�6�<�f=D��F�c=D�9�<��W0��f ����T��w�Ⱦ+ԟ���t�I�3�j���x   x   ;-���8�~$��$��8�5-��$���OE��z=��D}�5���ФȾ���_y	��v�=p&�ח/��T4��T4�ח/�;p&��v�ay	����ϤȾ/����D}��z=�VE�6���x   x   �?�c��־��y���?������ǽ�4���@��F}�c֟�O>¾��LZ�({������� �����'{�LZ�
��L>¾e֟��F}���@��4��ǽ����x   x   E�f��e�9��C�Z���D�ʽ�5��}=�D�t�|�m�̂Ҿ���x> �����D��D����}> ����ɂҾs�~�@�t��}=��5�B�ʽm���$�C�x   x   �TӼ����!UӼ�-��kE�@�����ǽNH���3��d�U���ﾤ�)��оyl߾h�3V�q�sl߾о/��𾤾P����d���3�XH���ǽF���skE��-�x   x   �ʫ��ʫ���μa-�|�C�򜉽��������]<$�oM��3w��􏾟A��(=��ۻ�=[��9[��ۻ�-=���A�����3w�}M�X<$�����x���윉���C��-��μx   x   ����ļ@[򼡟!���]��՗��J̽-����)��^P��(w�|̍�!�������J^��V���O^���������z̍��(w��^P���)�/���J̽�՗�_�]���!��Z�ļx   x   p ļ$�ؼ�����$��0V��U��|K���F�e-�Ծ-��J���e���{�첅�J͉�J͉�粅���{�ȑe��J�Ͼ-�j-��F轀K���U���0V���$������ؼR ļx   x   �E������N+��O�C��x����½`�뽽�9����1��?��I�]3L��I�"�?���1�7����j�뽲�½�w��R���O�Z+�O�����E�̱�x   x   ��!�|$�}�*�:7�`�J��g�9'��ۻ���^��aսm�Z���*��}��}��*�X��m�pս�^��л��G'���g�z�J�
7���*�7|$���!��� �Ć �x   x   r�]�mV���N���J��	L�*qT�Ƨd�|�?S�����YE��hJ��1�����1��[J��qE������2S��*|���d�5qT�w	L���J��N�VV�f�]�� c��)e�� c�x   x   5���A�� f���g�YeT��G��B�y�D���L�[�W�ic���l�j8r�b8r��l�ic�E�W���L��D��B�j�G�keT� �g�-f��@��9���{����;���;��b���x   x   7*̽�.��`��
����d�V�B���)��M�NQ�����#����N�����#����_Q�N�\�)�d�B���d���`���.��P*̽��ݽ���ƌ�����ݽx   x   .��k!�+�½��{���D�xC��B�Ƽ�詼x㙼����j㙼�詼9Ƽ�B�C���D��{�뢞�"�½t!�+��������%��%������x   x   ��)�p�f��c?���;��;�L��=��ż�*��D9��n�i���n�"9��*��>�ż>�H�L��;��]?��l��w���)�υ@���R��^��b�^���R�܅@�x   x   �@P���-���
�x�ԽА��#�W�h���ʩ�`f9�����B/��A/�����f9��ʩ�u����W�Ԑ����Խ��
���-��@P�R=p�E����!��J+��F+���!��D���?=p�x   x   �w��J��}��C｝%��";c�������8E�/���M�� /�eD������*;c��%���Cｭ}��J�w�V������{������/ǽ������{����X���x   x   *���\qe�.�1�8��m(����l����8���N���.���.�{��^���Ú���l�n(��1��1�1�aqe�&���()���8��?%Ծgc�����gc�<%Ծ�8��&)��x   x   �z���{���?���E���r��������8�Kٲ�8���������r�?������?��{��z���G���'۾���ޘ���
�c'���
�������'۾�G��x   x   T�������K�H�
g�����r���U���"L9��L9�|���
��r�����g�K�H�𡅾O�����ξ�.�u,	��m������$���$�����m�x,	��.���ξx   x   2K�������L��g����Թl���-©�F��©�����l�����g��L�����=K����ھB��	���%��}2��:��m=��:��}2���%��G����ھx   x   곾������H����,���?c������ż��żƐ��?c��,������H�����곾xᾊt��y�zO1���A��ZM��sS��sS��ZM���A�zO1��y��t�{�x   x   _M��t�����?�P��Y+����W��;�e,�;��W�N+��K����?�t���eM����Y	���!���8�<lL���[���e���h���e���[�;lL���8���!�Y	���x   x   ~���؉{���1�
N�%���e�L�t>�q>�l�L�-���N��1�ى{�w�����ھv���!��(;�R���d�%qr�_�y�c�y�'qr���d� R��(;���!�v���ھx   x   Ѐ���{e�Յ���Խ�A���D��)��D��A����Խυ��{e�׀��*�ξD���|���8�-R��h��*y�Q
��AꃿN
���*y��h�.R���8��|�G��&�ξx   x   H�����J����J���{��B��B��{��J������J�F����O��H7�I�vS1��oL�P�d�(,y��ڃ����������ڃ�(,y�P�d��oL�vS1�I�C7��O��x   x   �w�K�-�ߗ�l����d�ȻG���d�s���ۗ�J�-��w��2��'2۾2	�?�%��A���[�Cur����k���啉�k������Cur���[��A�?�%�2	�)2۾�2��x   x   �PP��"�J�½���jT��jT���G�½�"��PP�g����D���"���t��2��aM�A�e��y��샿9���8����샿�y�A�e��aM��2��t��"���D��h���x   x   ��)��7�n����g�jL��g�n���7轓�)��Qp�S��e3Ծ��������:�&|S�~�h���y�W���܃�X����y�{�h�&|S���:�������i3ԾY���Qp�x   x   O���A��}���J���J�}��A��J���@�]���(����s⾀���$��w=�k}S��e��yr�2y�2y��yr��e�n}S��w=���$�~��s�!���^�����@�x   x   YB̽�P��yO��7��O��P��dB̽����R��/��糺�p��h1���$��:�eM�)�[�"�d�h� �d�,�[�eM�ݭ:���$�g1�v��쳺��/����R����x   x   �ї�{-V�+�$+�S-V��ї�(޽y��2'^��:��ٽ���I����q�2��A�wL��R��R�wL��A�s�2����K���ٽ��:��,'^���>޽x   x   ��]�v�$������$���]�햠���齍�%�� b��;��y���cx���Ny�i�%�[1���8��2;���8�[1�l�%�Ly���ax⾁����;��� b���%����ۖ��x   x   g�!�������X�!��Ac�!T��*��ŝ%�y*^��2������:Ծe,��-8	���^����!���!�^����+8	�k,���:Ծ����2��o*^�ȝ%�)��3T���Ac�x   x   Y_򼖼ؼ�_�V� ��Le�.U�������(�R�3���A&���M���=۾yE���|�fc	�����yE��=۾�M��A&��4���2�R�����3U���Le�D� �x   x   �ļ�ļm��� ��Cc�����w޽z����@��]p�����=���\��S�ξ��ھ�%��%���ھV�ξ�\��=�������]p���@�p��o޽�����Cc�� ����x   x   s�ȼ[ ڼ��u�5�G{�ˬ��>�z�7RB� `n�B��C롾����;u��ʾW;ʾ;u������B롾!B��`n�8RB���>� ˬ��{�|�5����P ڼx   x   ��ټ���F��[=9�qr�����	н����.%��G�Pkh��`���現�՘�Xz��Sz���՘��現�`��Akh��G��.%����н����qr��=9�e������ټx   x   �y��~���#�9�@��Qj��Q��v���d߽�B�����U7��$L��l\�q�f�nZj�w�f�m\�x$L��U7�ƽ��B��d߽w��R���Qj�E�@���#��~��y�pM�x   x   ��5��+9��@��N���e���������M��0rս_����&
��,�$� ��%���%�� ��,��&
�^���'rսN��-���������e���N�)�@��+9���5��4���4�x   x   B�z��Qr��:j�i�e�I�g��r��A��rc��a{��񹴽��ŽW+Խwݽe��wݽI+Խ��Ž�[{��c���A���r�M�g�n�e��:j��Qr��z�ܳ���ၽ곀�x   x   ٯ��兟��>��q能L�r��>e�5�`��d��wo���}�_��;-2��(2��V[��y�}��wo���d�K�`��>e�a�r�^能�>��ۅ��߯��Ŷ��9���9���Ķ�x   x   7���Ͻ�洽'����3����`�6�E�8�4�g,�$U)�X�)�Z+�9,��Y+�C�)�+U)�f,�F�4��E���`��3��4����洽��ϽE��}���e�=���e��}��x   x   j��@���@߽]1���N���d�7�4���@��)�ּlƼ�f��'g��$lƼI�ּb����J�4��d��N��c1���@߽9��m��m*���6�=P=�5P=���6�h*�x   x   �4B��%�r,�QNսm`���Ro�V�+�����u����Q�yAB�7�Q� u��]����O�+��Ro�^`��ENսo,��%��4B��+\���p���}��/����}���p��+\�x   x   �=n�P�F����5��������u}�C7)�ftּg�����}�л��л���;g��etּZ7)��u}�����<������M�F��=n�`D��$v��i��F%��G%��i��!v��ZD��x   x   �.��2Ih��87�
���Ž0���
�)��@Ƽn�Q��лf���̓лC�Q��@Ƽ��)�,�����Ž
��87�.Ih��.��%��=���&TʾߺԾMؾٺԾ(Tʾ?���#��x   x   �֡�nN��oL����Խ(Ӌ��3+��5���B��oл�oл�	B�*6���3+�2Ӌ��Խ��nL�oN���֡�t���o�ھ��� ������� ���u�ھq���x   x   姳��ԏ��L\�C� ��Oݽ����+��4����Q�9��@�Q��4����+����rOݽ@� ��L\��ԏ�秳��׾�d��Mi�!��#�P� �#�"��Hi��d��)�׾x   x   U_��h�Q�f�E�%�s��9��4+�<ƼY��BY��&<Ƽ54+�G��r��M�%�W�f�c�L_����j�	� ��$+���5��;��;���5��$+�! �f�	���x   x   �ʾ�g��R;j�U�%�-Rݽ9Ջ���)�kּ#���^kּ��)�(Ջ�RݽZ�%�D;j��g���ʾ����8����)�"�<�.XK�)�T��X�.�T�)XK��<���)�=������x   x   ��̾�h��D�f�J� ��	Խ ���7)���󼥭�!7)� ����	ԽM� �E�f��h����̾f�������3���I���\��yj�	�q��q��yj���\���I��3����j���x   x   �ʾ;Ř�|R\�{�p�Ž�{}�8�+��y�2�+��{}�d�Žq�vR\�<Ř��ʾ������58�<_R��Vi�dM{��b���[���b��`M{��Vi�>_R�48�������x   x   d��Tُ�+L�

�;���QXo�%�4�*�4�LXo�A���
�9L�Uُ��c��&���u��@8�XDU���o�2���f���)��	)��h���1�����o�YDU�B8�s��$���x   x   }���FT���A7�p����g��4�d��E�>�d��g��x����A7�?T�������뾠���3��aR��o��ӄ��񎿠i��ȣ���i�����ӄ��o��aR��3������x   x   �ޡ�Vh�׭��[սeU����`���`�lU���[սխ��Vh��ޡ�3�׾;�	�l�)�}�I��Zi�����j�{�������~���h򎿳����Zi�~�I�j�)�9�	�:�׾x   x   �7��cG��6��=���8��;e��8���=���6�eG��7��
Ŀ�^p��l���<���\�+S{�����ek������b�����dk������*S{���\���<�l�_p��Ŀ�x   x   <Pn�r"%�VS߽×����r���r�����YS߽s"%�1Pn�����۾�p��,+�S`K�݁j�ef��f,���������������h,��ff��݁j�P`K��,+��p��۾���x   x   �FB� ��=���������g�����E�������FB��O��(
�������	6���T�֣q�3`��K-��4m��B���9m��J-��0`��ףq���T�	6����#��/
���O��x   x   ���н1L��Q�e�=�e�3L��н����A\�����~dʾ� �S-���;�	X�S�q�h��f�����������c���h��W�q�X���;�S-�� �udʾ⃘��A\�x   x   �4�ܗ��Oj���N�Oj�ᗟ��4��2*�%�p��x��c�ԾL ��� �+�;���T�=�j�XY{�����؄����[Y{�:�j���T�,�;��� �N �g�Ծ�x���p��2*�x   x   3Ƭ�umr���@���@�Qmr�0Ƭ������6�q�}��6��\aؾ2!�a/�|6�feK���\�|ci�J�o�M�o�|ci���\�ieK�~6�a/�1!�Qaؾ�6��t�}��6�����x   x   �{��?9�,�#��?9��{��޶�<x��h=��?���7��M�Ծ�� ����2+���<�?�I��kR�PU��kR�B�I���<�	2+������ �W�Ծ�7��~?���h=�2x��޶�x   x   N�5�&�����I�5��ƀ�'V�����5j=�.�}�`|��jʾC��%v�s���)��(3��!8��!8��(3���)�p�+v�I��jʾ\|��-�}�@j=� ��6V��ǀ�x   x   d���񼇈���4�����[W��%z��6�2�p�[������0۾�}��G�	���&��)�&���I�	��}��$۾��a���3�p�$�6�z�_W������~�4�x   x    ڼ#ڼ"\�)�4��ǀ�ⶽԥ��)9*�oK\��V���!��п�٬׾�%뾮���� �� ������%�֬׾п��!���V��mK\�$9*�ԥ��$ⶽ�ǀ�K�4�Q\�x   x   ��ؼ���k����G�����ܿ�����*��Y������������6HȾZu׾.�RF�9�Uu׾3HȾ������������Y��*����ܿ�������G�%�����x   x   %�� �?���bK�텽bF��轫����8�\�^�S���oْ�� �����ͯ��ͯ�
���� �vْ�L���V�^���8�����]F��텽�bK�^��'�F��x   x   ������S3���S�-��������ʽ
,��ƹ��M3���M�?e�\Gw�1l���g��4l��fGw�-e���M��M3�����+���ʽ����)�����S��S3���q���x   x   �G��NK�}�S��d���~�"���2����̽����
���ĺ*��o5�W;�^;��o5�ɺ*�����
�����̽�2������~��d���S��NK���G�$`F��_F�x   x   P���xۅ�?�����~��"��?ԇ��ѓ�9���������ͽ>���-�����ZM ������-�<�Ὀ�ͽ����F����ѓ�9ԇ�#����~�:���vۅ�*����:��8����:��x   x   Y����+��D}��3���̇��-���m�����򉽲В�"����̢�[���Q����̢�#����В�������m��-���̇���R}���+��c�����ʽRѽ`ѽ��ʽx   x   (������ɽ��C��^�?&c�t[R���J�?�I�o)L�M�N���O�,�N�B)L�L�I���J��[R�)&c��^�+�(��#�ɽ���'���.�w��*0�~���.�x   x   �*��j������̽x��`���NR��-��s������ٴ��J���������s�ӈ-�*NR�`���*x����̽����j�(�*���=�ںK��S��S�޺K���=�x   x   ��X�J�8����d��y��މ�F�J��h�'��Kx�����l������Bx��Ж��h�/�J�މ��y���d���Z�8���X���u��2��)������+����2����u�x   x   � ��i�^��03���
���ͽ1���)�I�F��h��QRx��gD�=hD�Sx�&i��J�C�I�4�����ͽ��
��03�f�^�� �����5橾�
���i���i���
��1橾���x   x   d���n偾W�M������ ���xL������f��RTD��E �BTD�2f�����TL������ ��P�M�j偾f���7뷾 Ͼ�4ᾆ�쾳��}�쾒4� Ͼ4뷾x   x   �t��+Œ���d��*��ڭ��!�N����ׄ��JD��ID�.�������N�뭢�3��*���d�+Œ��t���zվA��[�i\�����h\�[�K��zվx   x   P0Ⱦ�����#w�8S5�'���˚��֯O��~���_��$2x��_���~����O�њ�����4S5��#w�����P0ȾO��*�
�U���'�c0���2�e0���'�P�)�
�Z��x   x   *]׾�{Z���:��7 �����ޙN������Z���Z��������N������7 ��:��Z��铪� ]׾��]'�ܒ-��>��J��:Q��:Q��J��>�ߒ-�Y'���x   x   e��9����V��9�:�1���T���{L���~����L�I������<�:��V��8���p�ྺ[
��B$���<�'"R���b�F�m��_q�L�m���b�!"R���<��B$��[
�x   x   �/�F���\���V5��򽑙����I�-a�1a���I�������V5�"\��L����/侉O�JB+��wG��Ca���v��6��`O��_O���6����v��Ca��wG�KB+��O�x   x   �����+*w�K�*�ɲ�������J�r|-���J����²�B�*�"*w������]P��-�mM���j�$���ތ��|��*ŕ��|��ތ�%�����j�kM��-�]P�x   x   Tb׾�����d����m�ͽ�ችXIR�aIR��ችs�ͽ�����d�����Ob׾(^
�AD+��M��$n��C�����cB��������gB������C���$n��M�AD+�&^
�x   x   �7Ⱦ�˒�ʴM��
����������c����������
�ƴM��˒��7Ⱦ���\F$�{G�D�j��D���"��ܠ�9b��~���3b��ܠ��"���D��?�j�{G�`F$����x   x   �}���쁾><3�t�����_��_����t�;<3��쁾�}��\�ﾸ,�+�<��Ha�k�������ܠ�A㪿)��
)��D㪿�ܠ����l����Ha�)�<��,�`��x   x   X���%�^�@���̽.ȓ�,��6ȓ��̽?��'�^�X���s�վ��
��-�l)R���v�iጿ3E��Hd��*��ز�*��Gd��4E��hጿ��v�l)R��-���
�s�վx   x   ���8����O'��|Ї��Ї�A'������8�������������>���b��;��D����"������>+��;+�������"��D����;����b���>����������x   x   ��X�y��ʽ����$������ʽy���X�����%Ͼ�c���'���J�k�m� U���ʕ��#��cf��}檿if���#���ʕ�U��n�m���J���'��c��%Ͼ���x   x   Q�*����\�����~�{�~�c������V�*��u�t����F��f��0��FQ��lq��U��"���0H��	ᠿᠿ,H��%����U���lq��FQ��0��f��F�x�����u�x   x   ����?������`d������?�����g�=�1A��?����V�[�2�3HQ�}�m�>���䌿O��S(��Q���䌿>��z�m�6HQ�]�2�W���=��+A��`�=�x   x   x׿�녽��S���S�녽׿�'A���K�!���}��1��V�&0���J���b���v�Z���iJ��kJ��Z�����v���b���J�#0�U�)��}��&�����K�5A�x   x   '���;eK�u^3�GeK�%����˽��U:S����`~��M�쾣i�C�'��>�o1R��Ra��j�2n� �j��Ra�t1R��>�A�'��i�U��b~�����V:S����˽x   x   ��G���������G�<P��7ѽIF��;S�4���& ���L�ph��!�ġ-���<�e�G�hM�mM�h�G���<�¡-��!�rh��L�" ��8����;S�NF�*7ѽMP��x   x   ��}$�+���|F�ئ��v8ѽ9��Y�K�E������:.Ͼ����
��5��P$�8P+�0�-�6P+��P$��5��
����>.Ͼ����E��Y�K�%��w8ѽ�����|F�x   x   *��R�뼒��|F�ZQ���˽&E�V�=���u��'��@����վ� �y���h
�Q\�N\��h
�|��� 𾲓վE���'����u�U�=�+E��˽`Q���|F���x   x   �㼙���z���U�y��b�ϽQ��!:���l�(��⫾�ľ�<ھ	�����Ρ�������꾣<ھ �ľ⫾(����l��!:�Q�]�Ͻ�x����U��z����x   x   ���i
�G�(��Y�x���D_�������-"��J�-�s�����������j���������j�����������)�s��J��-"�����G_��y���B�Y�a�(�1i
�,��x   x   �k�$�(���?�2�c�$*��˯���ܽ�	�W�&��D�gb��{��ć����PA������ć�؟{�db��D�O�&��	���ܽ˯�#*��=�c�V�?�'�(�sk�А�x   x   mrU�&�Y���c��Nv�q��C �)G���s��(p���,��=�B�H��&O��&O�:�H��=���,�p�n���DG��< �q���Nv���c�V�Y��rU� T��T�x   x   9b��3m�����li��""���{���ƣ�Q���lν���z������>)������y������lνQ��hƣ��{��,"��pi�����9m��b���2�������2��x   x   ��Ͻ�A�������Zs���r��0:��UI��JE��c:��$����t��D��:���t��)���`:��VE��DI��=:���r��]s��۱�������A����Ͻ@�۽�g��g��۽x   x   H:�"���T�ܽ�-�������1��4X��o�s��n�@p�<�t�
�x���z��x���t�@p���n�y�s�2X���1�������-��X�ܽ���C:��l��k!��4$��k!��l�x   x   �:��"��	�5���7���9���s���N��7�+�*���$�;"��;"���$�Q�*�#�7���N��s��9���7��<���	��"��:���N���]���e���e���]���N�x   x   ��l���I�Ut&���� Lν�.����n���7���� ��eB���ټBἡ ������7���n��.��Lν���Kt&��I���l��Ņ���v�)���w����Ņ�x   x   q��bvs���D��V��������p�L�*�e��nl�����������l�����_�*��p������潿V���D�`vs�l������⸾�ƾ��̾��̾�ƾz⸾����x   x   
˫��	����a�l�,��N���ز���t�F�$��'�_���-��\���p'�R�$�a�t��ز��N��w�,���a��	��	˫��?ȾJL����7� ����2� ����HLᾭ?Ⱦx   x   S�ľ#n���z{���<����?S���x�b"� �ټU���)���D�ټp"��x�YS�������<��z{�!n��Y�ľ^辈���$����!!�#!�����$����^�x   x   �"ھ퐯�y�����H��������qz�"�H!�)\��7!��"�qz�����r��}�H�x��������"ھ&����,�(�2�6���?���B�ź?�2�6�(�(���+��x   x   ���T�����]O�<�{���e�x���$���������$�d�x�����F�iO����T��֜��C�í&��	=�=�O��E]�Kbd�Cbd��E]�D�O��	=���&��C�x   x   )���p뿾�.���	O�8��(V��M�t���*�����*�f�t�*V��,���	O��.��o뿾1���ܑ�V�2���M�^`e�x����N������
x�Y`e���M�W�2�ّ�x   x   9����쿾}��H�H����ݲ�p���7���7�p� ݲ����L�H�����쿾7���a���:�v�Y�o-v�0!��ߏ�Hz��Gz��ߏ�2!��k-v�r�Y��:�d��x   x    ���W��괇���<�hW���#��'�n���N�"�n��#��eW����<�䴇��W�� ��H��[ =���_��m��)�����44��rɤ�04�����+���m����_�V =�H��x   x   v��`���K�{���,���R3���s��s�D3������,�U�{�e���w�꾀��3�:���_��C���I��d���4 ����������8 ��`����I���C����_�5�:�~��x   x   �*ھ.u���a�_�,Vν�<���S���<��"Vν_��a�*u���*ھH�~�2�@�Y�Uo���J��S���V��u乿�ؼ�n乿�V��Y���J��So��?�Y�~�2�H�x   x   �ľ���A�D�4���@�� 3��3���@��4��?�D�����ľ�����&���M�43v����Z���X��S����¿�¿V���	X��Y������63v���M���&����x   x   �ի���s�ـ&��Ὓ����q��������؀&���s��ի��j�;���=�mhe�2%��ս��d#���湿&�¿��ſ&�¿�湿d#��ս��2%��lhe��=�;���j�x   x   ����I��	�P;��	x��x��C;���	��I����qMȾ���&�(� �O�Jx�I䏿-9�� ���\ܼ�n�¿k�¿Yܼ�$���-9��G䏿Ix� �O�%�(����sMȾx   x   ��l��#"���ܽ����n$��������ܽ�#"���l��Ħ�]ᾬ.��6��Q]�
�������Ϥ�O���1鹿���8鹿N����Ϥ�����
���Q]��6��.�]�zĦ�x   x   �:�����^į�-q��2q��kį������:�3Ӆ�󸾸�����V�?��od�}������I;���&���\���\���&��M;������{���od�T�?��������;Ӆ�x   x   ]K�xX���(���Xv��(��nX��^K�Y�N�����ƾd� ��$!���B�iqd����珿�������������������珿���lqd��B��$!�b� ��ƾ���W�N�x   x   ��Ͻn~���c���c�t~����Ͻ����]������̾���%!���?�V]��x��)��B$��<Q��>Q��A$���)���x�	V]���?��%!�����̾����]����x   x   �v���Y�[�?�	�Y��v���۽�!���e�󽜾[�̾$� �����6���O�Qqe�C>v��u��K���u��H>v�Tqe���O���6���(� �[�̾潜���e���!��۽x   x   ��U�}�(�e�(�̏U�oJ������L$�C�e����ƾ����3���(�1=�1�M���Y��_��_�Y�+�M�1=���(��3�|���ƾ��Q�e��L$����rJ��x   x   �}�Or
��}��'T�u���'��Y�!���]��!������pf�ْ�>��h�&�
�2�V�:��.=�S�:�	�2�k�&�@��Ԓ�qfᾬ����!����]�F�!�$��j����'T�x   x   q�����Ң�0'T��K����۽��ذN�م��̦��XȾ+y�e��gR�E��K��H��F��kR�_��,y辮XȾ�̦�م�ٰN����۽�K��J'T����x   x   _��j2��\Q!��^��.��_ܽ�&�s:F��\|�ؚ�	`��)�Ѿ���(c��}��v�����c�����2�Ѿ`��ؚ��\|�y:F��&�Sܽ�.���^�HQ!�m2��x   x   �%����2�.��c�Me���*̽���L-�w(X�(g���*���ث����g�Ǿ|;|;i�Ǿ����ث��*��(g���(X��L-���+̽Ne��$�c�>�.���A&��x   x   MA!�r�.��G��co�䄔��z��ɧ콯T�,L3��/T� �s������A������^������A������ �s��/T� L3��T�ħ��z��߄���co���G�}�.�!A!�M�x   x   �u^���c�XVo��a����������O�ͽ�0������'�'<���M�!�Z���a���a��Z���M�*'<��'�����0��a�ͽ���������a��^Vo���c�v^���\���\�x   x   {���P���u�������ؗ�tG��:��z�ɽd6�į�����V������ ���_���������u6�}�ɽ:��fG���ؗ������u���P��U���֠�>���֠�x   x   ��۽�̽�a��&����>�����;r��u馽~��>�����̽��ֽ�tܽ�tܽ�ֽ��̽;���~��`馽Dr��<����>������a���̽��۽{>�M��Y��d>�x   x   E�{�� �� �ͽ0(���i��F�=8���ƌ���|��J���5ݗ�X����|�������ƌ�>8��R�i��(��'�ͽ��y��>��"�-+��-�6+��"�x   x   WF�1-�J=����ܼɽ�ئ��0��M`x��d��Z��V�ͩU���U��V��Z��d�I`x��0���ئ��ɽ���J=�1-�hF�؏[��Nk�ܢs�ɢs��Nk�ڏ[�x   x   �6|��X��/3��y�佞f�����.vd��B���-�2{#�J] �,{#���-��B�9vd�����f��佗y��/3��X��6|�_W���9��V���\��W����9��eW��x   x   &��S���T�1�&����nڿ�o���j�Z���-��s�q�q��s���-���Z�p���|ڿ� ���)�&��T��S��#�Ry��:�ľulҾƭپϭپslҾ5�ľRy��x   x   �G����Yus�o	<���b�̽Cg���V��m#�l�k%��l��m#��V�0g��P�̽��{	<�Wus����G��v8վ<���5�$��Q ����5�9��o8վx   x   ��Ѿ����;z��U�M�H��g�ֽ)���G�U�xM ��i��i��M �7�U�'�����ֽT��R�M�8z��~�����Ѿav����݀���%��l+��l+���%�؀���_v��x   x   v�����-����Z�����Qܽ�ŗ��U�$k#�l�"k#��U��ŗ��Qܽt����Z��-����w�辌��� ���3�|�B��\L�P�O��\L�}�B���3��� ���x   x   xG��mlǾ����ȅa�����Rܽ/���O�V�z�-���-�C�V�����Rܽ���ׅa�����flǾnG��X��e�1�O�I�h�]��Ql��t�~t��Ql�n�]�L�I�d�1�X��x   x   ߬��d;�K��M�a�h����ֽ�h���Z��B� �Z��h����ֽa��C�a��K���d;��qu �:�>��[�h'u�Ƿ��)?������.?��ŷ��f'u��[�8�>�lu �x   x   t���e;s����Z����R�̽���_pd�gpd�����;�̽����Z�����e;t���%���F��ah�����Pڐ�hl���y���y��gl��Qڐ������ah���F��%�x   x   t��pǾR1����M�Ȏ�࿽����pUx�¹��"࿽Ȏ���M�K1��pǾq���%���I�.o�芉�����F[��(���.p��%���H[������ꊉ�)o���I��%�x   x   iM����Y���<�1���
l���/���/���k��6����<�[����oM��Ex ���F��o�����7/��H �����7���=������B ��4/�� ����o���F�Cx �x   x   ���ɫ���s�N�&�s��ܦ��쒽�ܦ�j�T�&���s�ɫ���՗���>��eh�����.0��5���2P��r�ȿZ̿j�ȿ3P��;���,0�������eh���>�ٗ�x   x   V�Ѿ���bT����2�ɽ�k���k��=�ɽ��aT����U�Ѿa���1���[�Ӻ��ʛ��r��iQ����˿_�ҿb�ҿ��˿eQ��p��͛��Ӻ����[���1�^�x   x   0S���\��"=3�^��c0������i0��W�� =3��\��2S������@� ���I�*0u��ސ�d_�������ȿ��ҿ`ֿ��ҿ�ȿ����e_���ސ�)0u���I�@� �����x   x   Κ�/X�J�Y�ͽ@D��PD��O�ͽJ�1X�Κ�Gվ@�+�3���]�a���r������"���Y̿,�ҿ)�ҿV̿&�������r��b�����]�*�3�C�Gվx   x   N|�%B-�Y��5����ۗ�'���_��B-�N|�'�����9��&�B�y^l��E�������v��q�����ȿ��˿��ȿp����v�������E��z^l�)�B�6����#���x   x   �0F�O��%t��L���R���1t��Q���0F��e���ľV@��%�[jL�[t�r�����������N����V��}V��K���������p���Vt�WjL��%�Y@��ľ�e��x   x   � �$̽ȃ���g������$̽� �M�[�=J����Ҿ���z+�z�O��t��G��/u���c��0��4���4���c��-u���G���t���O��z+�����Ҿ3J��R�[�x   x   Sܽcc��Vjo�Vjo�qc��eܽq�"��kk�Փ��-�پ`-��{+�mL�)cl�����}㐿ݡ��j7��k7��ޡ��|㐿����.cl�mL��{+�a-�3�پᓣ��kk�t�"�x   x   �,��n�c���G�h�c��,���`�A+���s�p����پ���_&�V�B�O�]��9u���������������������9u�G�]�X�B�e&������پp����s�;+��`�x   x   e�^��.��.���^���!��.�o�s�.���"�Ҿ�C�r��S�3��I��[�:sh��'o��'o�=sh���[��I�S�3�s���C��Ҿ9���|�s��.��!ｵx   x   �T!����T!���\��X���"ｧ +��pk��N��˰ľ����Ƚ �'�1��>���F�#�I���F��>�(�1�˽ �����ְľ�N���pk�� +��"ｏX����\�x   x   �8���8����%�\��𠽐d���"�&�[��k��󐱾�Rվ�����Ϣ�ʄ �� %�� %�̈́ �Ӣ�������Rվ��k��*�[���"��d���+�\���x   x   U����N�!��5b��i��������N�c���-�������9�۾�t�M�����v�
����C���t�D�۾|���-���a�����N���ג��i���5b�o�!�����x   x   ����Ĺ��0��h��R��6CԽ|����5��b��툾�ן�O���C�ž��Ѿ�׾�׾��ѾK�žF����ן��툾�b���5�v��NCԽ�R��?�h��0����A���x   x   ��!��x0���K�)�v�g���{ĽF��]��@�=���`�������q���0�������0��v��}������`�1�=�U��
F��{ĽW���$�v��K��x0���!�z�x   x   �b���h�K�v�˲���?��= ���a۽�[��F�
�3��qJ���]���k���r���r���k�~�]��qJ���3��F��[��a۽< ���?��߲��9�v���h��b�^�_�v�_�x   x   �P���=���t���7��(���j�����½��ܽ��������%���&��&.�Խ0��&.���&��%����������ܽd�½\���2����7���t���=���P�����l���x   x   �m��"Խ:aĽC��C���~���@^��'���˽�۽�C��<��/���(����<���C��۽�˽'��E^������F���9��CaĽ�"Խ�m��s�|������s�x   x   ���&��� ��zE۽	�½ZU��缧�_1���}���$ٳ�����8:�������س������Z1������IU���½xE۽
!��%������(���0�e�3���0��(�x   x   CjN�j5�3���H�N�ܽ���)���/���?��\��񍽏n��xn���q򍽴?���/���)����Z�ܽ�H�3���i5�WjN�6
d��s�r_|�[_|��s�9
d�x   x   ؛��@�b�ǭ=�/�����˽⧽�9���ˁ�k�s���l���j���l�r�s�{ˁ��9��⧽˽����/���=�O�b�؛��E���1��á��g���ġ���1��J��x   x   �����و��`���3����۽펭�5荽W�s��M]��XS��XS��M]�X�s�I荽���۽�����3���`��و������Ը�2e̾בھ{⾆�ґھ*e̾ ո�x   x   S�������H��RSJ����"뽦ó�L卽׎l��SS�XxK��SS���l�H卽�ó��"뽹�^SJ�H������K����8޾h���g�OA�W��JA��g�	h���8޾x   x   e۾�r������s�]�V�&�W���k���`���~j�RS��QS��~j��`���k��v��c�&�t�]�~����r��"e۾����v�!���,�+u2�,u2���,�q�!�����x   x   �X�rž�욾ek��.�k���v#���`���l�;G]�2�l��`���#��Z����.��dk��욾�rž�X�G���'�d;�XK��$U��X��$U�XK�d;���'�I�x   x   ����ѾB��r�r�֥0�Ǜ��Lm���卽��s���s�~卽6m�������0���r�M��	�Ѿ���:�pN9�3dR�\�g���v�������v�b�g�.dR�pN9�:�x   x   ����׾ے���r�.�Q���ų��獽ǁ��獽�ų�f���.��r�͒��	�׾����'�UG��ge�t:������瑿�M���瑿���s:���ge�PG��'�x   x   �
�S�׾E��sik�j�&��(뽞���8��8�������(�g�&�qik�S��Z�׾�
�!h,���O��s���-헿$"��j���i���#"��-헿�􉿥s���O�%h,�x   x   4���Ѿ��^�]�*�á۽�㧽|+���㧽ס۽-�j�]����Ѿ1��%i,���R��%z��*���H��������Ϻ�������H���*���%z���R�&i,�x   x   ���xž�A\J�F���	˽�)���)���	˽F��5\J���xž���'�)�O�E'z�]N���2��X%����ÿʿ	ʿ��ÿQ%���2��`N��K'z�/�O��'�x   x   �a�jz���	��u�3���������������������3��	��kz���a��>�G�s��,���3�����s�ɿ��ӿ��׿��ӿu�ɿ����3��,��s�G��>�x   x   p۾�ʟ�T�`�>9��ܽ�X���X��*�ܽ:9�S�`��ʟ��o۾e�U9�ne�����K���'����ɿsa׿��޿��޿wa׿��ɿ�'���K������ne�U9�`�x   x   a����㈾6�=�wR���½;�����½uR�5�=��㈾d���-���'�mR�?�����j�ÿ��ӿ�޿6A��޿��ӿj�ÿ���?��mR���'�-�x   x   �����b�΢�+V۽'���8���V۽֢���b����?H޾���-n;���g����>(���Ƿ�O"ʿ݅׿��޿��޿څ׿T"ʿ�Ƿ�:(�������g�+n;����?H޾x   x   ���|5��8�����1������9���{5����~举�z��V�!��K�zw�ݎ��׺��#ʿp�ӿ�e׿w�ӿ�#ʿ�ֺ�����zw��K�P�!��z��~举x   x   ��N�֬��tĽPA��OA���tĽܬ���N�%���w̾�r���,�)3U�~)��U�� ���(ʷ�n�ÿ?�ɿ9�ɿk�ÿ/ʷ�����U��w)�$3U���,��r��w̾%��x   x   ����<ԽɃ��d���˃���<Խ����$d�C����ھ�M�y�2��X�(+��𑿈+�������-������-�������+����.+��X�w�2��M��ھC���$d�x   x   ��\Q����v���v�oQ���㽌�(�ft�
����������2�6U�kw��������R��y;��y;��R���������qw��5U���2��������bt���(�x   x   Fh��K�h�9�K�6�h�1h�������0���|�7���t⾴O��,�%K�G�g�7D��{��� 4��W��4��~���7D��>�g�%K��,��O�p�)�����|���0����x   x   �7b�h�0���0��7b�rä�Y2��A�3�^�|�o�����ھAv���!��u;��vR��ze�Ls��7z��7z�Os��ze��vR��u;���!�=v�|�ھ}���l�|�K�3�Q2��fä�x   x   [�!���(�!���_�
���3��/�0��t��G���~̾��������'��_9��!G���O���R���O��!G��_9���'��������~̾�G���t�"�0��3��#
����_�x   x   ��������!�U�_�hĤ�����(��,d�S+����]T޾��%�8J��'��w,��w,��'�=J��$���gT޾{�P+���,d���(����iĤ�D�_�|!�x   x   �$ؼ�z����v`����c�@���R����X��� �ľ	?����{�y�C��y�
{����?���ľY�������R�3��sc����v`�����z�x   x   [m��	��.�4i��X��u�ؽ"a�U�:���i�"a���$�������7ܻ̾ؾB;߾8;߾�ؾ�7̾�����$��#a����i�R�:�a���ؽ�X��64i��.���	��m�x   x   ����.�t�K�z�uh���˽>��R["��OF��k�I��[���9�������Q�������9��[��I���k��OF�J["�C���˽]h��z�x�K��.������x   x   ?W`�zi�z��k��z���o����`������%���?�NSX���l���{�$���0�����{���l�gSX���?���%�����`�h���u���l���z�|i�ZW`���\���\�x   x   | ��]C���X������
۪�����k�ӽI��
��q��d+��38��}@�i[C��}@��38��d+��q��
�D��T�ӽ~���۪������X��zC��Z ��S���]���D���x   x   >���ؽl˽]��`}��9w����ƽ	ֽ{齍)����(������*�����)��{��
ֽ��ƽTw��d}��S��q˽Òؽ>�m2�#E��#E��d2�x   x   ����J��z�}D���ӽǡƽR���KĽ��˽S�ս�߽���P9���彀߽e�ս��˽�JĽd�����ƽ�ӽsD轧z��J����_�*�7�2�wW5�H�2�L�*�x   x   u�R�g�:�
C"�˲���<�սrCĽ���tt���>���2���;���;���2���>��ht��/���pCĽ1�ս ��ڲ�C"�Q�:���R���g��$w�\^�C^��$w���g�x   x   V�����i�2F�#�%�0�	��c��˽�n���ӯ�$Ϋ�����.s������+Ϋ��ӯ��n���˽�c�8�	��%�2F���i�X����ʖ���������䮾��������ʖ�x   x   {����L����j���?�]���~�ս�4��rʫ��ۣ�i���y����ۣ�jʫ�5����ս.��]���?���j��L��z���ك��>�Ͼ�޾�v��v徍޾5�Ͼー�x   x   �pľQ��}���B5X�N+�x�;�޽�&���w�������z�������&��.�޽x�N+�L5X�}���R���pľ��������	���	�����	�������x   x   �#�؀��+G����l�8����_��s/���l��죠�ߣ���l��f/��d�彗��'8���l�'G��Ѐ���#�z��M���$���/���5���5���/��$�U��z��x   x   �����̾`%��[�{��e@�l��V$��/�������٣�ך���/��f$�d���e@�N�{�Z%���̾�����j��+�@?�S9O���Y�U]���Y�S9O�@?��+��j�x   x   �l�,�ؾx���[���GDC�<��p���'���ɫ��ɫ��'��^��7��SDC�a�������&�ؾ�l���!�(n=�LW���l��|��n���n����|���l�FW�)n=���!�x   x   �j�B#߾Q>��8���h@����߽/6��ѯ�56���߽��h@�2���C>��>#߾�j�g�+���K���j��A���V���������������V���A���j���K�^�+�x   x   �w��$߾�����{�� 8��{�Đս�n���n����ս�{�� 8��{������$߾�w�p�0�Q�T���x��^���ԛ�hk��J��I��gk���ԛ��^����x�a�T�u�0�x   x   �l�.�ؾv)��^�l�T+����ݻ˽(���Ի˽���$T+�n�l�l)��#�ؾ�l�}�0�׾W����L֓������˳�����M-�������˳�����O֓����ʾW��0�x   x   �o�?%̾�L���>X�d�7l齪EĽ�EĽ3l�d��>X��L��F%̾�o�x�+�ܩT�a�����"���e��	Yɿ�5п�5пYɿ e��������e���T�v�+�x   x   �������`��B�?��
��ֽ����ֽ}
�R�?�_�����������!���K�q�x� ؓ�7���V]��I�Ͽ�ڿDC޿�ڿK�Ͽ_]��4���ؓ�p�x�{�K���!�x   x   �.�����k��%�����ƽ�ƽ���
�%��k�����.�6q��t=��j�sb������wg����Ͽ?$޿\��_��B$޿��Ͽug��囥�sb���j��t=�0q�x   x   �|ľ	W��PAF�7��O�ӽ�y��R�ӽ9��OAF�W���|ľ���+�hW��F���ٛ�[г�]ɿ�ڿ�忹�����ڿ]ɿ[г��ٛ��F��hW�+����x   x   l�����i�gQ"��V�Յ��煻��V�mQ"���i�i���n�⾄���J?�+�l��\���q�����W;п�G޿��忆���G޿];п���q���\��)�l��J?����l��x   x   򴆾�:�Q�����xઽ���X���:�����ȓ��+)��K	%�FO��|�1������4���<п�ڿ�(޿�ڿ�<п�4����4����|�FO�D	%�#)��ɓ��x   x   ��R��Z�]˽����픡�_˽�Z���R��ٖ�$�Ͼ�	��0�m�Y�w��U��@�����7aɿh�Ͽa�Ͽ3aɿ���C��R��	w��g�Y��0��	�*�Ͼ�ٖ�x   x   �����ؽ�h���s���h����ؽ�����g�R���3޾Ե�P�5��]��w��A���1u��Nճ��m��2e���m��Kճ�.u��>����w���]�M�5�ϵ�(޾L�����g�x   x   /^�X��=z�$z�(X��D^�}�*��Cw�N��������5�a�Y�+�|��`���ޛ�����EĪ�EĪ������ޛ��`��0�|�R�Y���5�����]���Cw�z�*�x   x   ���Q9i���K�19i����W��2�?�����C��·� 0��KO��l��K��i���������ߓ�i���K���l��KO�(0�÷�=������4���2�W�x   x   Yy`�%.�T%.�}y`�N����l���r5�������"޾��	��%�/R?�SW��j�!�x��$���$��&�x�x�j�YW�.R?��%���	��"޾�������r5��l��?���x   x   =���	������\�����n��9�2�Iw��ţ�*о_3�����&+��=���K�
�T�n�W� �T���K� �=�&+����]3��9о�ţ��Hw�*�2�	n��������\�x   x   �����w��b�\�����Z񽡾*���g���������	㾟���z�>"���+�)�0�'�0���+�C"��z�����	㾰��������g���*��Z����F�\�M��x   x   �WǼ? �
l��Z� ���������xS��t��Y禾�2ƾ�[㾮v��m��^��{�b��b���v���[�~2ƾY禾�t��xS����������Z�Al�J �x   x   �༤'� :(���e��ڽ��ʳ=���m����4a��3\���iоS<ݾu��k��Z<ݾ�iо*\��2a������m�ó=���+ڽ���e��9(��'�;�x   x   #[��/(�wH�p{z�3۠��4н�����'��M�3�s��<���$���|���M�������M���|��|$���<��A�s��M���'�����4н۠�c{z�!wH�0(�[�{��x   x   5�Y�gne��mz�rA��ߓ��<8ʽ	��4����0�q�L� g��}��u���������u���}� g�]�L���0�=��)	��68ʽۓ���A���mz�fne�S�Y���T���T�x   x   �����ڞ��ˠ��������yʽ���6���O�G-�+?�`qM���V���Y��V�qqM�?�D-�P�4������yʽ�������ˠ��ڞ�����/Ϡ��f��$Ϡ�x   x   ޸���ٽ=н�&ʽqʽ�Oҽ��὿���@�����4=!��)���.���.� �)�2=!����F��������὿Oҽqʽ�&ʽAн��ٽڸ����;��:�����x   x   ރ�����������ˠ�C���[��b������q�����y�������b���� \�6�ώ�罱���������Ѓ�u+)��O0���2��O0�c+)�x   x   �WS�i�=�+�'�¢�%���p�����e����{��P� �����T� ��{�����f�p��)��Т�)�'�Q�=��WS���f�X�t��|� �|�b�t���f�x   x   a����m�RxM�ߗ0�R?�8w�%V�����p��R�-�������,���R�k�𽅡�V��:w�Z?�ԗ0�FxM���m�a��"���ܱ�����iZ�����ܱ��'���x   x   �Ц����s�4�L��-�@�����s���N�ܘ�k�y�͘��N�s����N���-�3�L��s����Ц�����o#Ͼϸܾe��r��ɸܾf#Ͼ����x   x   tƾXK���*��Bg���>��.!���\� ������ُ������Z� ����.!���>�Hg��*��ZK��mƾz[�b���,<	���)F���7<	�Z���n[�x   x   �@��D��@��h�|�2[M��)�(�����/��� ��$������*���)�;[M�t�|�>���D���@㾌P�%��Ϥ$��r/�8%5�9%5��r/�ʤ$�-���P�x   x   �Z���Qо�h���f��ޞV���.��= �����U�ｯ���@ �Ɉ�ڞ.�֞V��f���h���Qо�Z���
�XC+��%?�9�N��(Y���\��(Y�8�N��%?�UC+��
�x   x   5��Q$ݾ :��3�����Y�ݟ.������ �"P�P�� ����ٟ.���Y�9���0:��M$ݾ/����"�L�=��.W���l��|�lr��er���|���l��.W�M�=���"�x   x   j��/���精���t�V���)�K
��v������v��S
���)�x�V�����精*��k���,�E9L�I k�!v��ő���Õ��A���Õ���!v��T k�?9L��,�x   x   4����S<��i��@`M��2!��z������2!�8`M�i��d<�����7��1��ZU�Osy�l����E���6���6���򦿸E��h���Jsy��ZU��1�x   x   &��n(ݾm��X}��?�����\��Gg�\������?�h}�m��c(ݾ"��%�1�A}X��y��qL���4�������ݽ����ݽ������4��tL���y��5}X�(�1�x   x   x��Xо*��yg��-��|����|��-�lg�-��Xо}��4�,�p]U�mz��U���Po���R���vʿ�nѿ�nѿ�vʿ�R��Lo��X���pz��v]U�1�,�x   x   �c��CM���1����L��G��z���^��z���G���L��1��CM���c����"�6>L��wy�MN��ip��cZ���ѿ��ۿ��߿��ۿ�ѿkZ��fp��JN���wy�0>L���"�x   x   CL�U����s���0���%��������0���s�U��@L�3�6�=�|'k�����8��/U��" ѿ��߿[�"[翲�߿ ѿ-U��8������'k�8�=�,�x   x   &ƾO���5�M���W�罩TҽW����6�M�M���&ƾ�W��K+��7W�	{���J�������zʿ�ܿ�\��K뿹\��ܿ�zʿ�����J��	{���7W��K+��W�x   x   �ݦ�F�m�8�'�����{ʽ�{ʽ���<�'�M�m��ݦ�fk�s��0?�Q�l��������>使^tѿ��߿]^�Z^翏�߿ctѿ@使�������P�l�0?�y��bk�x   x   �m����=�ݐ��6ʽT���6ʽ����=��m�����������$�O�)�|�W˕��������uѿ�ܿe�߿�ܿ�uѿ���!���[˕�)�|�O��$���������x   x   eoS�s�W1н�����\1нz�moS�s���q6Ͼ�G	��/��7Y��z���J��P����潿	ʿ�%ѿ�%ѿʿ�潿S����J���z���7Y��/��G	�v6Ͼt���x   x   ���ڽ�ܠ�@J���ܠ��ڽ���f��â��ܾ� �45�B�\��{��i͕����������[��]b���[����������g͕��{��N�\�45�� �u�ܾ�â��f�x   x   s�����z�w�z�
𞽋�佴B)�mu�ͯ��J��,T�:55��:Y�>�|�웎�P���>���x���x���>��P��𛎿B�|�~:Y�555�/T�R��ۯ��iu��B)�x   x   ����F�e��H�'�e�}������_i0��|��o�������1�/��O�9�l�M����č�?V��^���9V���č�M���0�l��O�9�/�����㾇o���|�\i0����x   x   �Z�1D(�hD(��Z�D꠽����2�r�|������ܾ-K	�x�$��7?��AW��3k���y�ς��ւ����y��3k��AW��7?�v�$�'K	���ܾ�����|���2���3꠽x   x   q��2��p��U������|k0�!u��Ǣ�/=Ͼ����H���T+�8�=�PKL��lU�̍X��lU�PKL�9�=��T+�F������>=Ͼ�Ǣ�u�ik0���*����U�x   x   �'��'����U��꠽���jF)�(�f�;���1���w㾎_���7�"�3�,���1���1�9�,�;�"����_�w�)���7���.�f�|F)����꠽�U����x   x   .�����˼�P��P����� �߽� ���P�<��j���v!ž?f�T���}��m�����r��t��[���Hf�q!žk���<����P�� ���߽�����P�Q���˼x   x   uy˼�*� �*O_�����fٽWw��>���o�`o��L2�����h�Ҿ��߾Զ�ɶ���߾o�Ҿ���J2��ao����o���>�Sw�)fٽ����<O_�� ��*�y˼x   x   @�< ��sC�n�y��񢽌ս]�	���-���T���|��c��졾���pݶ�Ф��oݶ����졾�c����|���T���-�b�	��սu�k�y��sC�I �d@�X��x   x   [ P��7_�T�y�H�������սO<��q�\�=���\�k�x��@���Ð��6���6���Ð��@��w�x��\�a�=��q�R<���ս���H��=�y��7_�w P��*I��*I�x   x   N����蜽�⢽)���������ݽ�� �z��-�]�C�n�X���h��s�)w��s���h�f�X�]�C��-�z��� ���ݽ����#����⢽�蜽4���>�����=��x   x   ��߽nGٽRս8�ս@�ݽ���B��$5��#���3���B�r}M��IS��IS�z}M���B���3��#�5�A�����J�ݽ.�սWսfGٽ��߽���̞�ɞ�~��x   x   ��@b��	�u/�� �_��\�	� ��s����+���5��<�-�>��<���5�Ĕ+�h����f�	�Y��u� �o/�)�	�Ab���B�$��~*���,��~*�6�$�x   x   ��P���>���-��`�n��-����Q ��!�w@)�&�/�K�3�F�3�)�/�{@)��!�Y �����-�r��`���-���>���P��Sa�L�m�
�t���t�T�m��Sa�x   x   u)���o���T�:�=��
-��#����!��e%�,�*��o.���/��o.�0�*��e%��!����#��
-�1�=���T�,�o�x)�������~������(������~������x   x   Ө���\����|��l\���C�>�3���+�6=)��*���,�y�.�~�.���,��*�?=)���+�G�3���C��l\�µ|��\��Ѩ��jR���Xʾ��־S�ݾ^�ݾ��־�XʾrR��x   x   q	ž����R���x�n�X�+�B�{�5���/��n.�G�.�[�.�H�.��n.���/�v�5�$�B�f�X��x��R�����k	ž<�߾N��o���?�Kp��?�x��N��3�߾x   x   pL��u��%ڡ�)3���h��pM���<��3��/���.���.� �/��3���<��pM�
�h�/3��&ڡ��u��uL�A������� �DD+��0��0�AD+��� ����A��x   x   w�����Ҿ笮�/����ss��=S���>�ܯ3��o.���,��o.�ݯ3���>��=S��ss�(���ݬ����Ҿ{����/�K;(��3;�~]J��-T���W��-T�|]J��3;�I;(��/�x   x   �t�I�߾�˶��)��%w��>S���<���/�!�*��*���/��<��>S�*w��)���˶�E�߾�t�7� ��:�ES���g�Dw�h3�\3�Bw���g�@S��:�:� �x   x   )���������*���vs�stM��5�u@)�h%�z@)��5�vtM��vs��*��Г����*���*���H���f��܀�G���+������0���D����܀���f���H��*�x   x   `��s���Ͷ�渐���h���B���+�]!�\!���+���B���h�⸐��Ͷ�z��b��ê/�R���t��	���;��]����6���6��\����;���	����t�R�ƪ/�x   x   ��w�߾L���q7��5�X���3� ��J#�&����3�5�X�w7��C���n�߾��ӫ/��*U�6p|�ፑ����2)���N���z���N��3)�����㍑�0p|�{*U�ի/�x   x   8x�_�ҾLࡾ�x���C�#�������#���C���x�Pࡾd�Ҿ;x��*��R��q|�F͓��D��۹�/�ƿ�Ϳ�Ϳ2�ƿ۹��D��H͓��q|��R�
�*�x   x   ى��d~��ZZ��y\�?-��4���	��4�?-� y\�UZ��c~��։��!� ���H�hu������E��Gݼ�~gͿ>%ؿ�ۿ6%ؿ�gͿNݼ��E������gu���H�&� �x   x   �W�p'���|��=���!�������=��|�u'���W�6���:���f�������ݹ��hͿ�ۿWf�Zf��ۿ�hͿ�ݹ��������f�²:�6�x   x   !žg��E�T�m��� �a��� �m�H�T�g�� ž����C(�jS��ဿ~@���-��6�ƿ9(ؿ�g�8N��g�8(ؿ6�ƿ�-��~@���ဿjS��C(����x   x   �����o�X�-�u:���ݽ��ݽm:�Z�-��o������߾��W>;�:�g�����Ʋ���T����Ϳ��ۿ�i㿊i㿭�ۿ��Ϳ�T��ò������9�g�W>;�!���߾x   x   E6����>�#�	���ս}���{�ս(�	�v�>�I6��eb��@a��!�+jJ�X(w������>�������Ϳ@+ؿ��ۿG+ؿ��Ϳ�����>������Y(w�.jJ�!�=a��fb��x   x   ;�P�^s��ս[���U����սcs�?�P�Λ��Ukʾ���@Q+�]<T��C�|$���?��rW��j�ƿ�nͿ�nͿf�ƿxW���?��y$���C�Y<T�CQ+����Xkʾћ��x   x   ���cٽ���_R��
����cٽ���na�a����־@L���0��W�^E�¶��'����2�� 乿"弿乿�2��$�������cE��W���0�=L��־[����na�x   x   �߽����,�y��y�����4�߽9�$���m�i���äݾ~���0�/?T�E-w�C����E������M���M������E��G���I-w�#?T���0�~�ʤݾt�����m�>�$�x   x   ����W_���C��W_�󵚽���*��t��=��6�ݾN��T+�poJ���g��怿���|���֓�x�������怿��g�toJ��T+�	N�2�ݾ|=���t��*���x   x   #P�8 �T �2#P��8��x���,�t�t�t���)�־��+!��E;��S���f��u��|�%�|��u���f��S��E;�)!�	��$�־������t� �,�p���8��x   x   QV�pB�'V�}NI�#7��A��ڙ*���m�4����qʾ}j����L(�J�:�.I�&R��:U�R�0I�K�:�	L(����j���qʾ0�����m�ƙ*�;��37��{NI�x   x   K�˼��˼� �#MI��8����C�$��ta�����*j���྽���>��� �u�*���/���/�x�*��� ��>������#j�������ta�T�$���8��MI�� �x   x   Qh���L����
�D�����0ٽ�/��{L�z��������.¾�O߾�i�����������������i���O߾�.¾����y����{L��/�ٽ�����D����L��x   x   
@���ܼ�B���X�M����Uؽ���h�?�yDq��r��̎��<¾��Ծ��
�� �辄⾊�Ծ�;¾ˎ���r���Dq�a�?�����UؽQ�����X��B�3�ܼ(@��x   x   ���9���>���y������۽���+�4��]��̓�����*�&[���ؾ�j����ؾ�)[��(������̓�ܸ]�-�4������۽�����y���>��9���*��x   x   ymD�uX�k�y��╽{��y��3��-��[O�q������
Q��8.��C.��Q�������q��[O��-��3�y�"{���╽d�y�uX��mD�&&;�&;�x   x   �k�����I���s��mjӽ߱��]��>,���G�I�b�{�����@��H^���@�����{�L�b���G��>,�]�ϱ��ijӽ�s��O�������k��������������x   x   �ؽQ9ؽ{�۽�i�g����	����N�0�cnG��O]��1p�~���������'~��1p��O]�hnG�J�0������	�x����i�|�۽F9ؽ�ؽ�۽�ܽ�ܽ�۽x   x   $�0t�ژ�+(��U�/��8})��:�8_M�m!_��m��\w��z��\w��m�t!_�6_M��:�>})�*���U�((���0t�%����	�!��c#��!����x   x   �^L��r?��|4���-�4,�-�0�e�:�glH�ƥW���e�$�p� �v�!�v�)�p���e�ǥW�flH�`�:�.�0� 4,���-��|4�vr?��^L���X���b�%h�
%h�üb��X�x   x   ���m&q�Y�]��HO�ӾG�GfG�[M�N�W�0�c�E�n�7@v�e�x�0@v�I�n�"�c�N�W�[M�GfG�оG��HO�O�]�v&q� ����������3����ӟ�3����������x   x   �碾Da������p�w�b�}F]��_���e��n��\v�+�z�2�z��\v��n���e��_�}F]�y�b���p�ￃ�Ea���碾�|��,¾�%;gӾnӾ�%;,¾�|��x   x   X¾�{����������]{�d(p�U�m���p�A@v���z�ޟ|���z�?@v���p�L�m�`(p�[{����������{��R¾�Xپ���j- �H��>��C��o- ���Xپx   x   �7߾�'¾F⨾����+��~��Xw�r�v�g�x���z���z�j�x�r�v��Xw�'~�.������H⨾�'¾�7߾������h�
�#�n�(�q�(�	�#�h�������x   x   �P���Ծ/K���E���9������+�z���v�uBv�z_v�zBv���v�0�z������9���E��+K���Ծ�P��"Q��m"���3���A���J�#N���J���A���3��m"�$Q�x   x   E��=�ɾ�b#���W��m����[w�.�p��n��n�)�p��[w�m����W��j#��ɾ�8�A��P���n4���J��[^��l��?t��?t��l��[^�~�J��n4�R��x   x   i��������s$��B;���~�i�m�3�e��c�6�e�r�m��~�B;��q$��ޱ�����k���]&��fB��*^��kw�����~��3ʎ�~�������kw��*^��fB��]&�x   x   ����o˾��H��~��R/p�x#_���W���W�n#_�N/p����H��{˾��辍��X+��CK� �k������������k"��j"���������������k��CK��X+�x   x   &��x
��O�������{�O]��bM��rH��bM�O]��{������O��q
�#���Y+�yNN��5s��ߋ�i��w㩿����������x㩿k���ߋ��5s�sNN��Y+�x   x   �����Ծ�訾���I�b��oG��:���:��oG�H�b�����訾��Ծ����`&�<FK�Y7s�A��ԃ���H��ť���7ſ�7ſǥ���H��҃��B��]7s�?FK��`&�x   x   Z���0¾����k�p�R�G�g�0�փ)�m�0�O�G�y�p������0¾Z��&��vkB�m�k�nዿ℡��0���ſ-QϿ��ҿ'QϿ�ſ�0��ᄡ�lዿk�k�ukB�*��x   x   C߾܅���ȃ��VO�U?,�o��k��[?,��VO�ȃ������B߾fW�:u4��1^� ���y���,K��ſ��ҿS$ڿV$ڿ��ҿſ+K��{��� ����1^�9u4�cW�x   x   �$¾�k����]�Y�-��_���	��_�`�-���]��k���$¾A����u"�d�J�uw������穿����TϿ�%ڿ��ݿ�%ڿTϿ�����穿����uw�e�J��u"�@���x   x   �����;q�^�4�~4�U���t���{4�[�4��;q�����%hپ��+�3��f^��慿H朿���=ſT�ҿj'ڿg'ڿR�ҿ=ſ���F朿�慿�f^�*�3���#hپx   x   ӱ��I�?�����~彌wӽ�~彧��E�?�ֱ��L�������r��A���l�e����)�������>ſ�VϿ@�ҿ�VϿ�>ſ�����)��g�����l��A��r����J���x   x   .vL����<�۽|���w���I�۽���/vL�鐎�S>¾@8 ���#��K�`Ot��Ҏ�+�����������ſ�ſ��������+���Ҏ�\Ot��K���#�B8 �U>¾퐎�x   x   -�Vؽ�"��&�"��Vؽ!-���X������:;u��s�(��2N��Pt�K���}霿�쩿NQ��G8��RQ���쩿z霿J����Pt��2N�s�(�s���:;������X�x   x   ^ٽ�Ú���y���y��Ú�qٽ6��9�b��ŝ��Ӿr����(�i
K�G�l�$ꅿ���Ј����������ψ�����&ꅿJ�l�`
K���(�r���Ӿ�ŝ�8�b�>��x   x   Q�����X�՟>���X�D���%:۽7�!��Dh��矾2Ӿ����#���A��m^��~w�����苿����苿����~w��m^��A���#���1Ӿ{矾�Dh�0�!�):۽x   x   �D��O��O��D�ћ���ܽ�|#��Eh��ǝ�>;S; ��w���3�5K��<^��l��Fs��Fs��l��<^�:K���3��w�O; �>;�ǝ��Eh��|#��ܽ͛��x   x   ���ܼ{��H;�'ʐ�z�ܽy�!�}�b�ҵ���C¾�����W}"��~4�)wB��SK�{]N��SK�,wB��~4�X}"�������C¾ѵ��y�b�g�!�|�ܽ.ʐ��H;�x   x   �T���T������F;�"����:۽O��XY�+���쒳��qپ����r_����l&��f+��f+� l&����n_������qپ撳�*���RY�\��;۽����F;����x   x   )����b���켿a9�[����ѽ&���^G����������}���_۾�J������	�����	�����J���_۾�}�����������^G�'����ѽ[���a9�����b��x   x   �V��b�ɼ����S�V���K�ؽ�{�AA�N�s�9$��0�����ľ��׾�W�c\�\\쾦W征�׾��ľ0���9$��R�s�AA��{�H�ؽZ�����S�$����ɼ�V��x   x   ��켗��c�;���}����~�彣1�1�>��Rj��a��q���ɲ�����	ʾ�;�	ʾ����ɲ�q���a���Rj�1�>��1�t�������}�F�;����g��ajܼx   x   nG9��wS���}�0���|ǽ������}KA��ag�<���M��"���~��${��+{��{�����P��;����ag�KA��������ǽ�����}�xS��G9�1�,��,�x   x   hF��o������8ǽ�/�&��[i*��J��<l�������������������������������<l��J�Wi*�"��u/�Aǽ���j���XF���@���c��A��x   x   �ѽ��ؽ��彘�������#�B=��eZ�W�x��֊��(��+$��4ा2ा2$���(���֊�V�x��eZ�D=��#�����������ؽ�ѽ:�ν1�ͽ,�ͽ%�νx   x   ����j��#�#x�@c*��=���T���o�������朾��������朾��������o��T��=�6c*�#x��#��j��������>�����x   x   �DG��*A���>�v>A�z~J�4aZ��o��E���ِ���q���쨾�쨾#q��"���ِ��E���o�9aZ��~J�|>A�~�>��*A��DG��N���T�p�X�k�X���T��N�x   x   Z���ƭs�l=j�SRg��2l���x�m����ِ������i����������i�������ِ�p�����x��2l�PRg�i=j�˭s�Z����,���ގ��x��f���x���ގ��,��x   x   ������V����������ӊ�Q�����j���Ҭ�C氾H氾�Ҭ�j��	��R����ӊ��������V����������������"`��(-ž,-ž&`����������x   x   �i������Hd��>��)��
&��b圾�q�������氾�Ų��氾�����q��]圾	&��,��<��Fd�������i��F�оed��u���}��l��� �fd�C�оx   x   J۾w�ľ����%���㗠�"��3���:��簾�簾�=3���"��䗠�#�������v�ľ�J۾�A��R����ĭ�8�;�ŭ���T���A��x   x   �4����׾���� �����ޤ���2慨����Gլ�Ź��1慨���ޤ�������������׾�4��|
�̆�n�)�'6��C>��A��C>�'6�l�)�Ά�~
�x   x   ����F�L�ɾ�s��e|���ߤ����^t��mm��lm��Zt������ߤ�e|���s��Q�ɾ~F徖��0>�4�+�,�?��'Q�1^���d���d�0^��'Q�*�?�1�+�/>�x   x   s�	�<L�o;�t�������$���蜾2��#���3���蜾�$�������t��e;=L�v�	�c� ��K9�'R���h��Z{������˅������Z{���h�,R��K9�a� �x   x   ���M���ɾV��ܛ���*��;����ސ��ސ�9����*��ޛ��V����ɾ�M���wp%���A��H_���{����R��헿헿S�������{��H_���A�yp%�x   x   -�	��J徴���c������Yي�ǅ��J��ǅ�[ي����e��������J�+�	�{q%�,�D��.f�(Ã�s��SU���^���)��^��RU��u��*Ã��.f�)�D�{q%�x   x   ݷ���׾{ò���������x���o���o��x��������~ò���׾߷�]� �&�A�Q0f�nӅ�ս��r:������a¸�f¸�«��p:��Խ��nӅ�T0f�'�A�[� �x   x   2>��P�ľ�l��:����@l��mZ�1�T��mZ��@l�@����l��M�ľ0>���B��P9�!M_��ă�վ�����G���x8¿%�ſr8¿H������Ծ���ă�M_��P9��B�x   x   �U۾ۮ��"_��Ibg�N�J�/'=�,'=�U�J�Ebg�_��ܮ���U۾�"
���+��$R��{�W���<��������ſ�S̿�S̿��ſ�����<��X���{��$R���+��"
�x   x   tv������Oj��MA��o*��(#��o*��MA��Oj����tv���O�������?���h����Y��e���);¿\U̿��Ͽ\U̿(;¿e����Y������h���?�����O��x   x   ����^�s� �>�@��������<���>�`�s�����j�о���"�)�a2Q�.f{�"��%d��uǸ�G�ſ�V̿�V̿E�ſxǸ�&d��"��,f{�`2Q�!�)����l�оx   x   ䷀�?A��3�����A콽����3�?A�䷀���Nv�3���26� ^�z���&���s0���ȸ��=¿Єſ�=¿�ȸ�o0��'���z���^��26�2��Qv���x   x   �[G�E|����+ǽ�+ǽ��?|��[G�;��&����񾥹�'Q>���d��Ӆ�+���mf����������������qf��-����Ӆ���d�"Q>������&���;��x   x   ���T�ؽJ�����R��N�ؽ�����N���s��z���m�b%A��d�4���"���]��^B�����`B���]��"��2����d�h%A�o�v����s�����N�x   x   ��ѽl��� ~�	 ~�c�����ѽa���	U�6���]BžO0��^�xS>�-^��l{����*���ŗ��ŗ�*������l{�0^�rS>�\�L0��bBž7����	U�m��x   x   �^����S��<�ÙS��^���νߙ�%�X��-��fCž6���N��76��8Q���h�#�{��˃�"ۅ��˃�(�{���h��8Q�76�P��;���hCž�-��)�X�י��νx   x   �i9�k��F���i9��Y��ν�U��X������v���!�?����)���?��.R�CY_�T>f�Y>f�DY_��.R���?���)�?���!�v�������X��U�ν�Y��x   x   b�켾�ɼ��켄-�`|���νz���U�I�w���&}���M��0�+��Z9�J�A���D�I�A��Z9�1�+�N����'}�{���L񎾮U�i���ν]|��s-�x   x   Tk��lk��Q�ܼ��,�JX��;�ν=����N�>��"���оmZ��m)
�UK�R� ��|%��|%�R� �XK�i)
�qZ��	�о��>����N�F��N�ν<X����,���ܼx   x   �m�����Sܼ��0�D����c̽	���8C�*�|��˜��i���ؾc������'
����a��ؾ�i���˜�&�|��8C����c̽8����0�Sܼ
���x   x   U�������LW���R�:h��`�ܽ��	�E��y�#×�����ɾ|�ݾ��W��T����|�ݾ��ɾ�� ×��y��E���O�ܽ=h����R�iW�򼻼X���x   x   ~8ܼ�O�U�=�9;�������h��!�!���M���|�\����Z��wA����о��ھV�ݾ��ھ��оsA���Z��`�����|���M��!��h��ǈ��D;��+�=��O�&8ܼ�,ɼx   x   H�0�9�R��6���P��,�ܽj���2��\��S���3��#N������˾�WѾ�WѾ�˾���%N���3���S���\��2�m��5�ܽ�P���6��c�R�\�0��t ��t �x   x   򝉽�Y���~����ܽ<^��{&��K�'~s�bŎ�������:þ�@̾�ZϾ�@̾�:þ�����_Ŏ�'~s��K��{&�4^���ܽ�~��Y��ᝉ��y��)y�z�x   x   nI̽��ܽ�X����Ly&�l�E��	j�D��5n��ӓ������l�̾��Ҿ��Ҿp�̾����ϓ��4n��H���	j�h�E�Qy&����X����ܽxI̽��½Ӿ�Ӿ���½x   x   qu�.����!�"�2�K��j�S��q;�����)���rϾ<�ؾ��۾8�ؾ�rϾ+�� ��r;�� S���j�K�#�2���!�*��uu����3���U�6�����x   x   P"C�e�E�EM��\�
xs����
;���׮�����xҾ��޾{征徼�޾�xҾ����׮�;�����xs��\�@M�i�E�V"C��C�?�E�\G�\G�>�E��C�x   x   >j|��xy���|��M�������l�����;����Ӿ�>�~��8�v���>��Ӿ<�������l�������M����|��xy�6j|��|���"���凾w눾�凾�"���|��x   x   ��������~��e-�������������yҾ�?��.��������.?⾗yҾ����������l-���~���������L����}���+"��,"������ ���H�x   x   �X��{
���P��
H����y���tϾפ޾y��ؙ������ؙ��t��٤޾tϾy�����H���P��{
���X��RpǾk Ծ-߾:��aT�2��-߾n ԾPpǾx   x   �ؾ��ɾ�7��%���8þL�̾�ؾ�徏�9���6��������ؾL�̾�8þ%���7����ɾ�ؾ@�����e�e��<�<�f��d����=��x   x   
�𾩋ݾ]�о�˾@̾��Ҿ��۾T�)�뾲2�,��R���۾��Ҿ@̾�˾^�о��ݾ���f��^�x��/$(���.�B_1���.�0$(�u���^��f�x   x   ��·뾆xھ8TѾg[Ͼ
�Ҿ��ؾ̨޾�D⾷D�ʨ޾��ؾ�Ҿc[Ͼ;TѾ�xھɇ����%�a�!�΅2�DA�MPL��<R��<R�MPL�DA�υ2�^�!��%�x   x   z�Y��q�ݾ�UѾ�B̾�̾yϾ�ҾĻӾ�ҾyϾ�̾�B̾�UѾk�ݾY��}�&8���.��C��XW��cg�1�q�D�u�5�q��cg��XW��C���.�%8�x   x    
����K{ھ�˾�=þ`���d!����������f!��_����=þ�˾N{ھ��� 
����]�6��P�ݯh�0~���&\��$\��
��0~�ٯh��P�]�6����x   x   2�B�뾱�о4�����2����"��ா�"��1������3����о@��1����3�9�ߍV���s��^���O��x������x���O���^����s�ލV�2�9����x   x   9���ݾ.?���O�����u��pC��rC��u������O��2?����ݾ9�;���6�;�V���w�κ��4���+ˣ��@���@��.ˣ�2���̺����w�>�V���6�
;�x   x   B����ɾ�Y��;6���ʎ�V��[��T���ʎ�@6���Y����ɾB��^*���.��P��s��������QB���ޱ�)ݴ��ޱ�RB���������
�s��P���.�^*�x   x   �ؾ��ڈ���V��_�s��j��j�c�s��V��ֈ�����ؾ�l���!�"�C�ٵh�5a��B���xC��Qܴ�{��~��Sܴ�vC��B���6a��ڵh�"�C���!��l�x   x   $e��������|��\�)K���E�*K��\���|�����!e�����mf�Í2��`W�V8~��S���Σ�J᱿���Y6�����I᱿�Σ��S��V8~��`W�č2�of����x   x   �Ȝ���y�^�M���2�o�&�s�&���2�\�M���y��Ȝ��~Ǿ��������MA�Vng�^��)}��*E���ി
��
���ി,E��*}��^��Ung��MA���������~Ǿx   x   �|��E��!�i���i�h���!��E���|�����m1Ծ��.(�!\L���q��b������VF���㱿ി�㱿TF�������b����q�$\L��.(��q1Ծ����x   x   �8C�h���u����ܽ��ܽ�u��_���8C�u��������@߾q��/�VJR���u��c��2���ѣ�H��H���ѣ�5���c����u�UJR�/�r���@߾����y���x   x   Ԉ���ܽB��� c��G�����ܽՈ��	D�2���������HH��l1��KR���q�����W��V������X����W�������q��KR��l1�JH���澻���2���	D�x   x   �h̽wq���H���H��gq���h̽��sF�F����5��4k�I�	/��_L��sg�H@~�^f����������^f��D@~��sg��_L�	/�I�-k��5��F���tF���x   x   ߵ����R��>���R�ٵ��1ý|��jwG�p���}6����澞���2(�dSA�yhW���h���s�.�w���s���h�{hW�_SA��2(������澀6��j���owG�r��*ýx   x   d�0��g��g�a�0�8��k�&k��wG���������D߾R�g��g�2���C�&#P�u�V�x�V�'#P���C�g�2�i��T��D߾��������wG�&k�v�D��x   x   �bܼ�ػ�Acܼ�� �|Wy���G��=F�f3��{����6ԾI����k���!���.���6�٠9���6���.���!��k�B����6Ծ~���i3��?F�:����aWy��� �x   x   �%��Pɼ+� ���hýN��D
D�������>�Ǿ����q�1�&C�����%C�1��q����A�Ǿ������<
D�R��uý��I� �1Qɼx   x   b8Y��ꅼ݅Ӽ&�,��ㇽ qʽ)O���A���z���:e���7׾d4�6�����m�	����6��^4�7׾@e����~�z���A�0O�)qʽ�ㇽ1�,�:�Ӽ�ꅼx   x   v߅����,��AQX�4T��aA�I^�{�N�M^������&?��][Ӿ%辇���,���)�������)�d[Ӿ!?������Q^����N�I^�LA�;T��NQX�O������e߅�x   x   �lӼq��בF���G2ǽ��U}2��Lc��۬��/��f6־|p�c]���g]�{p�`6־/��ެ��󋾷Lc�Q}2���N2ǽ����F�\���lӼ8��x   x   0�,�hBX�3���Z�������m#���O����难�ʹ��̾u]�\��������Z��y]��̾�ʹ��难����O��m#������Z��>���BX�5�,�������x   x    ԇ��G��*ǽy���̽��GG�W5v��Ք��a��t�ȾHq߾�TQ��i �UQ���Hq߾s�Ⱦ�a���Ք�U5v��GG�ƽ�z���*ǽ�G��ԇ�Йr�"0i�ݙr�x   x   [ʽ�/潢���i#��EG���r�!i���a����Ⱦ��2��W*�}+�~+�W*�/���ᾰ�Ⱦ�a��#i����r��EG��i#�����/�[ʽ._���f���f��_��x   x   �@�tR��t2��O�w2v��h����ɾ���A��CX�Ώ�]��̏�EX��A�����ɾ򬾰h��w2v��O��t2�qR��@�>��TA�	� �SA�D��x   x   I�A��vN�Bc������Ӕ�!a���ɾ;��b� �@+���+
�-
���?+�c� �;�� ɾ a���Ӕ�����Bc��vN�N�A��:��G7��6��6��G7��:�x   x   ��z��U��틾q暾�`��݌Ⱦ٣�Ϗ �i��������!������i��Џ �գ���Ⱦ�`��m暾틾�U����z��v��v���w�k�x���w��v��v�x   x   x���1��������ʴ���Ⱦa��'D��c,�w���� �EV%�DV%��� �x��a,�*D��a����Ⱦ�ʴ�����/���v���፜��N���D��v��w���D���N��܍��x   x   �W��/5�� ��[�̾�q߾�
��;Z������0W%���'�0W%������;Z��
���q߾Y�̾���/5���W���Ͼ�2�ž�;̾Ѿ�Ҿ�Ѿ�;̾2�ž�Ͼ�x   x   �)׾xQӾ�0־\��,����,�t	!�*X%�+X%�w	!�,�����,��\��0־xQӾ�)׾p྿�뾿���� ��:��:�� ��������o�x   x   ]&����k�L���T���.�3���|��f� �x���1���.��T��H���k���\&�F3��c��	�����K)��
 �J)������a��L3��x   x   ���:���2Z���� �y/�w����������y��y/� ����9Z�8�����������7$�y�/��8�Ϗ=�͏=�߾8�|�/��7$������x   x   ���@���������(X��
/��]��0�^���0��]�	/�,X��������?������&U��#�+04��D�UEQ��Z�]��Z�QEQ��D�-04��#�&U�x   x   �	�ۆ��M]�ג�%���uM��'� �'� �xM�����$�Ւ�O]�܆���	� ��aV+��?�p�S���e��bs� �z���z��bs��e�n�S��?�aV+�!��x   x   ��������q�-c�Fz߾2��ڮ���ٮ�/��Hz߾-c��q������������-���E�j^�M�t������≿����≿����N�t�m^���E���-���x   x   ѿ�N�9־��̾��Ⱦ�Ⱦ�ɾ�ɾ�Ⱦ��Ⱦ��̾"9־N�Ͽ��W��X+�:�E�t�a�@�|�E>��'��Η�Η�)��D>��=�|�t�a�;�E��X+��W�x   x   �/� [Ӿ����Դ��k���l�������l���k���Դ����[Ӿ�/����#�ī?�J^��|��|��L��q������q��M��|���|�I^�ī?��#���x   x   �4׾>@��x���`��ޔ��s���s���ޔ�]�x���C@���4׾�>������54���S��t�@��T������.��0�����R���@���t���S��54�����>��x   x   -d��瞞�/���Lʀ�Gv�c�r�Gv�Mʀ�/���螞�)d���&�p���>$��D�|�e�Ń���t��T����K��T���t����Ń�|�e��D��>$�n���&�x   x   EÛ�Ka��DWc���O�6XG�4XG���O�FWc�Ka��DÛ�޾�R�뾁���/��NQ�Als�牿җ����{���y������җ�牿Als��NQ���/���P��޾�x   x   1�z�c�N�Ǉ2�{#�&��{#�ɇ2�a�N�1�z�����9�ž���������8��Z���z�W�� ӗ�3v�����7v��ӗ�V����z��Z���8��������=�ž����x   x   ��A��e����������e���A���v�s^��`M̾ � ��4���=��"]��z��艿��W���U�������艿�z��"]���=��4�!� �YM̾x^����v�x   x   �S�qO��Dǽ1q���Dǽ�O��S�S�:�[�v��U��x1Ѿ�E�� ���=�xZ��ps�Yȃ�}D��A���~D��[ȃ��ps�tZ���=�� ��E�}1Ѿ�U��N�v�R�:�x   x   YzʽLa��������9a��Yzʽ����_7��x�..����Ҿ.F�6���8�wSQ�*�e���t���|���|���t�&�e�zSQ���8�
6�-F���Ҿ2.���x��_7����x   x   
쇽?hX�t�F�_hX�쇽�}���T��36�ݧx��.���2Ѿ�� ������/��D���S�A^��a�>^� �S��D���/������ ��2Ѿ�.��ͧx��36��T��}��x   x   u-�v��=��n-���r�=���b� �z36�x��V���O̾G����D$��<4�R�?�X�E�Y�E�T�?��<4�D$� �L����O̾�V��
x��36�]� �O����r�x   x   �Ӽ����B�Ӽ+���Yi������S�%_7���v��_��$�že��>��Î�ʮ#��`+�;.��`+�Ȯ#�Ŏ�=��^��(�ž�_����v�&_7��S������Yi�&��x   x   �􅼆�3�����!�r��x��*��P�:���v�՜���྾-+ྏE������]������]�����E��.+ྑ྾Ԝ���v�L�:�&���x��(�r����f3��x   x   ��U�q턼�Լep/�f��|�ͽ�Z��&D�A�}������ּ��Dھ4�����%
�5L��%
����.���Dھ�ּ�����<�}��&D��Z���ͽL��bp/���Լo턼x   x   wℼY������f�W��������(�PL]�Z���A穾��Ǿ��)��y������x��.����~�Ǿ=穾\���SL]���(����e���f�������Jℼx   x   *�Լ���ZW��d��[߽����I�5���������nھ/Q�?��ž	����Ⱦ	�=��+Q�oھ	������3����I����Z߽�d���ZW�
��"�Լ�o��x   x   &^/��f��a����׽U��� @��v�{
��䗸�R�׾�d����S�� ��S�����d��S�׾㗸�y
���v�� @�[����׽�a���f�^/������x   x   =�������T߽���o3=��q�[Җ������/پ�`����
�&������K����'����
��`���/پ����\Җ�"�q�j3=�����T߽����9���$l��_��$l�x   x   ��ͽt���k��F@�B�q�<K��M����j۾C�����"���'��,��,��'� �����F���j۾M���9K��F�q�H@�n��r�����ͽ����%8��88������x   x   AO���(�J�I��v��і�c���SjܾHU�����+$���0� 9���;� 9���0��+$����IU�Ujܾc����і��v�H�I���(�DO��#�8u��.u��#�x   x   ]D��A]�빀�	�������k۾�U�pA���'��m7�x�B���H���H�v�B��m7���'�pA��U��k۾����	��빀��A]�^D���3�Č*��W&��W&�ʌ*���3�x   x   ��}�}���C���𖸾�0پ[�������'�2�9���G���P�|�S���P���G�0�9���'����\���0پ햸�C���������}���m��ge��ja�J`��ja��ge���m�x   x   e���"᩾��_�׾_c������-$��o7���G���S�+Z�(Z���S���G��o7��-$����^c��a�׾��᩾b���h���&#��]��W��W��]��)#��d���x   x   Jͼ���Ǿ_ھ/f����
�:���0���B���P�tZ�B0]�tZ���P���B��0�9����
�/f��[ھ��ǾOͼ��D���e�������^G������f�����D��x   x   7;ھ���jP�t�l��d�'��9�-�H�1�S��Z��Z�6�S�,�H��9�d�'�m��u�mP󾲧�4;ھ��ؾ�ܾX|�$��#��%��#��W|�ܾ��ؾx   x   $����������T��t�,���;�i�H���P���S�|�P�i�H���;�u�,�T����������'���9���
���9��B	����~(�����B	��9��
���9��x   x   ���&���	���	Q���,� !9�7�B���G���G�:�B�!9���,�Q����	�%�����I�i��M����Ċ$��(��(�Ċ$���O��j���H�x   x   1"
���������O����'���0�vu7���9�ru7���0���'�P����������5"
�]��FR�·$��]0��e:��+A���C��+A��e:��]0�·$�FR�^��x   x   �I�u����	����;��1��4$���'���'�4$�1��<�������	�v���I�p��ӟ �GL/��>��L�-}W��J]��J]�-}W��L��>�FL/�ӟ �p��x   x   �#
��������4�
������I� ����3�
���������#
�c���!#��4�}�G��Z��.i��1s�W�v��1s�.i��Z�~�G��4��!#�c��x   x   ��(���Y�9q��p������]��]����p��8q���Y�'����$��� �E�4��K��a�~�t�����ꆅ�ꆅ������t��a��K�E�4�� �$��x   x   ��� ���ھ��׾�>پ�z۾zܾ�z۾�>پ��׾�ھ�⾶��dM�:V��O/��G�Ma�I�x��օ�f ��{Q��e ���օ�I�x�Na��G��O/�:V�bM�x   x   �Fھ��Ǿ��� ��������ȷ��ȷ�������������Ǿ�FھE������$��>�=Z���t��ׅ��j�����������j���ׅ���t�<Z��>��$���� E��x   x   ڼ�������
ߖ�fX��	ߖ��������ڼ���ؾ�� ��d0���L��4i�(���F"�������`������F"��(����4i���L��d0� �����ؾx   x   f���ꩋ��ŀ�_2v�àq�àq�\2v� ƀ�멋�c����R���ܾ�A���$n:���W��9s�t���TT����������TT��u����9s���W�#n:����A��ܾ�R��x   x   ��}��X]�$�I�,3@�\G=�43@� �I��X]���}���$ ��݌��K	�R�$�y5A��T]���v�J���$��gm��$��J�����v��T]�y5A�S�$��K	����% ����x   x   �.D�[�(�@��x��p��<��`�(��.D�nn��1������]�澪��E((�̚C�3V]��<s�����ۅ�ۅ������<s�4V]�̚C�E((����\�澻����1��yn�x   x   �b������s߽�ؽ�s߽�����b�&�3�сe�Xl��"������53�	)(�n7A��W��9i���t�K�x���t��9i��W�n7A�	)(�23����(���Wl����e�'�3�x   x   ]�ͽ����y���y��񺬽R�ͽ�6�2�*�a�a��f��qY��b�龸��x�$��q:��L�LZ�a�a�LZ��L��q:�y�$����a��iY���f��l�a�8�*��6�x   x   �%���*f��}W��*f��%��³�M��n&��d`��f������1�澧M	� �Ii0�!�>���G�:K���G�!�>�Ki0� ��M	�0�����f���d`�n&�O��³�x   x   +�/����e���/�ZPl�fS���:�6m&�h�a�@l������9���C�����$�	V/��4��4�	V/���$����C�=�ᾓ���=l��o�a�:m&��:�xS��zPl�x   x   �ռ����ռa��A_��P�����}�*�Me� 1��� ���ܾ�����Z��� ��(#��� ��Z������ܾ� ��1��Ge�|�*�ɔ��P���@_�e��x   x   I��� ���Y������gEl�5����1���3��n�5
���Q��!�ؾcG���O�_��������^���O�gG��!�ؾ�Q��3
���n���3��1�8����El��������x   x   �d��Ս���ἁ49����d׽Q}���K�����⊣�H�þ٣�{v��9)	�������9)	�wv��գ�I�þ劣�������K�Q}�k׽���t49����Ս�x   x   �ʍ���ȼI[ ���|�v'�������9�E#s�HV�������H۾�-��4��7���|��|�5��5���-���H۾����DV��I#s���9�����'��	�|�A[ ��ȼ�ʍ�x   x   ���>V �j1q��Բ�����-�/�"�h����_T��Ǩھ�F��p���J� ���	"����J�o���F��ƨھgT�����!�h�/�/������Բ�l1q�EV �����¼x   x   �$9��|��Ҳ�����N�+�ipd�-)�����!޾(���O���!���+�=\1�>\1���+���!��O�*��޾����-)��jpd�T�+�����zҲ� �|��$9�������x   x   ?��/ ��������+�-Uc�F��N%��[�⾨f�Ǝ��2,�J�9�S�B�۔E�Q�B�K�9��2,�Î��f�^��Q%��E��'Uc���+�����2 ��D���m���\���m�x   x   �
׽�����/�nod�J���۹��w�\�	�h� ���5��G��wS���Y���Y��wS��G���5�g� �Y�	��w��۹�M��pod�~�/�����
׽����ނ�������x   x   �t��9�X�h��(���%���x徉�)2$��4<��<Q�!�a���k�^wo���k� �a��<Q��4<�+2$����x��%���(��Y�h��9��t�� �S���r߽H��� �x   x   &�K�>s�󛔾������e�	��2$�R�>�g�V�
�j��Vy��i���i���Vy��j�h�V�N�>��2$�f�	��⾊���򛔾:s�"�K�^41��� �Ia�Ea��� �Y41�x   x   ����ZS���S���޾dh�� ��6<���V�8n�d>��c	�����c	��c>��8n���V��6<�~� �bh��޾�S��\S������L�i�_�W���M���J���M�[�W�P�i�x   x   @���(�����ھ �����f�5�,@Q���j�&?��������������(?����j�)@Q�g�5��������ھ ���>���MF��P������������S��IF��x   x   ��þhG۾LI���R��6,��G�!�a�[y��
������������
��
[y�$�a��G��6,��R�II��mG۾��þK	��B���o���{;��wߦ�;��p���@���P	��x   x   #���-������!��9��~S�N�k��l��s��������u���l��J�k��~S��9��!�����-�����.վ��ξ!;R�;6Iξ5IξP�;!;��ξ�.վx   x   �r�����M�<,���B���Y��o��m�����@�������m���o���Y���B�<,��M����r���|�5ﾧ�����K��ne��J��������5��|�x   x   5(	������*c1�v�E��Y�;�k��_y�KB��MB���_y�6�k��Y�z�E�+c1������1(	��b�������|�&��
�
�&��x��������b�x   x   ���y��"�Ld1�
�B���S���a��j��@n��j�ğa���S��B�Ld1��"�z���|�����e��k�$�έ(�8Z*�ͭ(�$��k��e����~�x   x   e�r��œ��,���9�2G�
HQ���V���V�
HQ�/G���9��,�Ɠ�s��_���>���( ��H*��*4���;�E@�E@���;��*4��H*��( �=����x   x   �������Q��!�x=,�}�5�T@<���>�V@<�|�5�w=,��!��Q������� �����C%��2��?��BK�R�R�!�U�U�R��BK��?��2��C%������x   x   �+	��	�7���Y������ �E=$�A=$��� �����Y�8���	��+	�D�8���D%� T5�
�E��U��`���f���f��`��U��E��S5��D%�:��D�x   x   �|��d9���V����q��	��#��	�q����V��_9���|��
g�]���+ �`�2�U�E���X���g��q��qu�$�q���g���X�X�E�a�2��+ �^��g�x   x   9�⾘T۾�ھ�"޾���k��h�徣��#޾�ھ�T۾4�������j�kM*���?��U�S�g�B�u��=}��=}�A�u�V�g��U���?�lM*��j�����x   x   !�þ�����b��?����6��+��6��@����b������*�þ�;վGB�F���q�a04� HK�t�`�I�q�,?}�����,?}�H�q�u�`� HK�_04��q�F��CBﾩ;վx   x   �����`�������7��9��=��7�������`�����������ξ�����$�; <�"�R���f�rvu��@}��@}�tvu���f�!�R�= <��$���	���ξ���x   x   r����6s���h���d��nc� �d���h��6s�t����S��zƬ�40;������i�(��M@�@�U��f�3�q���u�-�q��f�C�U��M@�h�(�������50;uƬ��S��x   x   z�K�m�9�_�/���+���+�Z�/�t�9�z�K�B�i����SШ���;�#��=��c*��N@�[�R�4�`���g���g�7�`�W�R��N@��c*�>��#����;TШ����D�i�x   x   ���������������������IJ1�ָW�����J��7Zξ�w����ķ(��<�1LK�V"U�ЇX�Q"U�1LK��<�ķ(����w��7Zξ�J�����͸W�LJ1�x   x   �+׽l>����`>���+׽R� �v!���M�� ��料eZξ�$������$�(44� �?�F�F�#�?�'44��$�����$��fZξ料� ����M�z!�K� �x   x   �%���}�IZq��}��%��b������t���J�? ���J���;�����
��t��Q*��2��Z5��2��Q*��t��
�����ߠ;�J��@ ����J��t����a��x   x   QI9��u ��u �>I9���m�������߽Js�I�M�K��JϨ�0;\�����bm��/ �J%�J%��/ �dm����Z��0;KϨ�K��K�M�Is���߽�����m�x   x   ���ȼ%�v�Ƥ\�t�����罠!�(�W���Ĭ�'�ξB����1������!��1�����B�(�ξĬ���$�W��!����j�����\��x   x   �፼�፼O�¼��1�m�^	��� ��A1���i��N��B���7վD��bf���:��7����df�H��7վB���N����i��A1��� �\	��j�m���,�¼x   x    �����l����J�I ���V�""�_sY���������iо�8�/���.�5M�Z��8M��.�/���8��iо�������YsY��!"��V�I ���J�������x   x   ����㼽&5�����w�ս���46P��G��'֫�wѾ;���y��t��ջ#��(��(�һ#�q��|��E���mѾ֫��G��=6P�ǯ�v�ս�����&5�u����x   x   ����f"5����!bνL�C�L������r���1־_���Í�)�$�72�ŷ:��=�÷:�"72�)�$����_����1־�r������B�L�L�#bν���v"5����_	ּx   x   ��J������`νL��}K��4���P��}�ܾ����̒1�C�B��MO��U��U��MO�?�B�ђ1�����u�ܾ�P���4���}K�P��`ν����p�J���!���!�x   x   �����սK��}K������X��]��
���$�L�=���S�`Od��n�m�r��n�`Od���S�J�=���$��
�^��X�������}K�K���ս�����w�"b���w�x   x    M���v�L��4��UY��W������*�wG���a�?w��3���,���,���3��Cw���a�wG���*����V�UY���4��l�L��� M���������������x   x   �"��3P������Q���⾚��3�,�t�L��j�P���ӽ���#���R���#��ѽ��N����j�w�L�0�,�������Q�������3P��"���)���׽#����x   x   �mY��F���s�� �ܾ��
���*���L�D:n��^�������囿Έ��Έ���囿�����^��>:n���L���*���
��ܾ�s���F���mY�>3�|��&��&�|�>3�x   x   -��<֫�84־{����$�FzG���j��_���������踧�A.��縧���������_����j�CzG���$�}��E4־=֫�+��|�k���N�п>���9�ֿ>���N�~�k�x   x   ���Ѿ���Ϣ���=���a�����K��������2��J9��K9���2������K���������a� �=�Т�����Ѿ��� ��E܄��v��m���m��v�G܄�� ��x   x   �hоu���j��*�1��S�<w�*����蛿򺧿Z:��^˱�Z:��򺧿�蛿+���:w��S�,�1�i��z����hо����ڤ�𨚾�o�� ړ� p��祥��ڤ����x   x   s9�4��E�$�]�B��Wd�o8��(������Z1��j;��i;��Z1������(��q8���Wd�W�B�B�$�5��k9��w־�ž�߻�����1���1������߻�
�ž�w־x   x   \��q���=2�zVO�T�n�w2��X�����������5����������X��w2��M�n�|VO��=2�q��\��:/��z���ܾJ�پ�پ��ؾ�پP�پ�ܾt��9/��x   x   1� �#��:���U�e�r�L3���)���뛿���������뛿�)��M3��l�r���U��:��#�1��r�����������"����������� �������������r�x   x   �P���(�y�=���U�T�n��:���Č�����d"�������Č��:��M�n���U�{�=���(��P�pO��
��
�C/�p,�_����]��v,�C/��
��
�sO�x   x   �����(�K�:�pZO��]d�&w������e���e�������%w��]d�sZO�I�:���(�������e��*���!:��"�~�$�~�$��"� :����*��e���x   x   �R�R�#�dB2���B�,�S��a���j��Gn���j��a�,�S���B�dB2�P�#��R����5��_��;�-g'�$/��]4�E6��]4�%/�)g'�<�b��4�����x   x   �4�{����$�@�1���=�ʅG���L���L�ʅG���=�>�1���$����4�GR��g�^����!�v�,��l7���?�XD�XD���?��l7�v�,���!�`���g�IR�x   x   �����+�����%���*�r�,���*��%���2�������Vw���
�}-�P���,�NR:�u�E�{}M�1P��}M�r�E�LR:���,�P�{-���
�Uw�x   x   bF�P������/����
���������
�6�����J���^F�:��N���O
�߸�rj'�o7���E���P��V���V���P���E�o7�rj'���P
�K����:��x   x   wоe-Ѿ�E־2�ܾ��V���/�ܾ�E־c-Ѿwо��־¯�p���4�;?��/�@�?��M�:�V�էY�:�V��M�A�?��/�8?��4�r��Ư���־x   x   ��w嫾9����c��l��	l���c��5����嫾��]��v�žV�ܾ����2��"�Wc4��\D��4P�s�V�w�V��4P��\D�Wc4��"��2����R�ܾt�žg��x   x   �'��U�������D�������D������U���'��s.��B褾����پ��������$��K6��]D�T�M�'�P�L�M��]D��K6���$���������پ��:褾n.��x   x   ��Y��LP��L�ėK�ȗK��L��LP���Y�`�k�$鄾z���"���پ3�����6�$��d4���?���E���E��?��d4�4�$���5����پ"������(鄾X�k�x   x   �1"�)��`�%%�#`�#���1"��S3���N�۞v�k}��`@��6
پ����j��["�p/�'s7��W:� s7�o/�b"�i������6
پ_@��l}��Ӟv���N��S3�x   x   �o�Qֽ��νs�νZֽ�o��&�x��(�>���m�	瓾@���پ���#4�xA��m'�>�,�A�,��m'�vA� 4�����پ@��瓾��m�)�>�u���&�x   x   �2��R����'��L����2��j��I���7��9���m�|��� ����پ?���5�����i�!������5�H����پ� ��|����m��9��7�F��k��x   x   ��J��E5��E5���J�Yx����:"׽�5���>�'�v�b����껾H�ܾ�
���
��.��������.��
��
��<�ܾ 뻾i���(�v���>�|5�M"׽���Vx�x   x   ����?�`����"�Cb��	�����H����N��ㄾ�⤾�ž��������
��g����g���
��������ž�⤾�ㄾ��N�E������	��Cb��"�x   x   �Ơ��Ơ��*ּ�"��w������G3�S�k�&��|
��|־82���s�HO�������GO��s�82��|־~
��&��I�k�(G3������*�w�e"��*ּx   x   �~������J���b���"���81�U�l��d��T��h|⾱������&�+})��&�������j|�]���d��I�l��81�"�����b�K�#���x   x   ơ��S���_P���E��ǂ-�{]l������ þ�Z�������.�X�9���?���?�V�9�
�.�������{Z�� þ�����]l�ɂ-�)�����`_P������x   x   "A��[P�����z�p�,��qn�p��m�ʾ���������,��A�F�P��Z�?&^��Z�L�P��A���,��������i�ʾ
p���qn�{�,��z�*����[P�:A����x   x   �b�+���y��i,�rJp�S����Ҿ������N;�<XT��i��w��d��d��w��i�AXT��N;��������Ҿ\���dJp��i,��y�!���b��W2��W2�x   x   �쭽r��N�,��Jp�L좾<־#S��'�ءG��e�2�����lb����mb�����1���e�ݡG��'�S�<־L좾�Jp�W�,�w��쭽�?��o�o��?��x   x   �����-��rn�U���	=־��	� -,�p�O�N�r��H���N������U���U������N���H��H�r�q�O�-,���	�=־V����rn���-�����½b���a���ɟ½x   x   e61�
^l��q��ҾxT��-,�k�R�*�y�j��M^��Y���Of���	��Pf��W���M^��j��*�y�f�R��-,�}T�Ҿ�q��^l�^61�00	�N�VIսN�00	�x   x   �l������ʾ6����'���O���y�Ȍ���,��z���S��	�ÿ
�ÿ�S��z���,��ǌ����y���O���'�0����ʾ ����l��A:��k� � ��k��A:�x   x   e���þ�������?�G���r��k���-���-��%Ŀb�̿��Ͽ_�̿%Ŀ�-���-���k����r�>�G���������þe��i�s�KuK���4��o-���4�PuK�i�s�x   x   	���_����uT;���e��K��=a��M|��[Ŀ(�Ͽ(�տ*�տ)�ϿYĿL|��>a���K����e�sT;�����_���
㙾���;
g��aY��aY�7
g���� 㙾x   x   �⾧��	�,�`T���S������W����̿u�տ� ٿu�տ��̿W������S����`T��,���� ��f����������􆾑����������n���x   x   �����&A��i��
��ᑟ��k����ÿ��Ͽ��տ��տ��Ͽ��ÿ�k��⑟��
��zi��&A�����x!ݾ����
���+I��즟�馟�+I�����}���}!ݾx   x   A��H�.�=�P��w�'i���\������ÿ[�̿��Ͽ_�̿�ÿ����\��%i���w�F�P�H�.�>������X2߾P!;X�¾�׽�I^���׽�`�¾W!;S2߾����x   x   k�7:���Z��r�}����]���m���Z��ĿĿ�Z���m���]�������r���Z�4:�k��
����Q��xྵ�ܾS*۾X*۾��ܾ�xྟQ����
�x   x   �&�@�?��3^�Yt��j��Ԕ��ű��΁��g4��́��Ʊ��Ք���j��Wt��3^�B�?�
�&��-��$w �<����A�������������A��;���!w �2���x   x   [�)���?���Z���w�	���W��/g���4���4��1g���W������w���Z���?�W�)����{9�T��b�������
���������
����e��Q��v9����x   x   ;�&��:���P��i�����Q��s�����	s���Q������i���P��:�>�&����T��{n�0W����|y�Jx�Օ�Px�|y����2W�}n�U�����x   x   ���.�E.A��iT�l�e���r��z��z���r�l�e��iT�A.A��.����`;�ko�)���=�w����!�^�$�W�$���!�|���=�&��lo�a;��x   x   "��x��$�,��_;�N�G���O���R���O�H�G��_;�,�,�v�� ����
�͉���Y��>�,����&��",�U.��",���&�+���>�Y���̉���
�x   x   �%����������'��<,��<,��'����������%�����+��k{ ����|��x��	�&���.�:�2�6�2���.�
�&�v��|�����n{ �'������x   x   ^��vq��������.a�'
�5a��������zq�c���.ݾe>߾\� �����G}���!��$,�F�2��d5�F�2��$,���!�H}�������\�l>߾�.ݾx   x   ���Fþ�ʾq$Ҿ�S־�S־m$Ҿ�ʾOþ������������-;��ྻL���
��|�J�$�U.�-�2�1�2�U.�F�$��|���
��L����ྡ-;��������x   x   �s��9��� ���$����������0���3����s���𙾪��۰����¾4�ܾ���S�� ����$�<&,���.�6&,���$�%��P�����2�ܾ�¾ް�������x   x   �
m�tzl�Őn�Cjp�Xjp���n�fzl��
m���s�Q��t(���U��y佾47۾�������}���!���&���&���!��}�������57۾x佾�U��v(��T����s�x   x   ;M1�ԙ-�	�,��,��,�љ-�DM1�-X:�\�K�� g�� ��	����j���6۾U�����
��~�����������~���
�K����6۾�j������ ��� g�e�K�3X:�x   x   A�����}��^�ｯ��A���B	�j~���4�vY�9�����1㽾3�ܾ�L�������hA�kA�������L��6�ܾ3㽾���;��vY���4�a~��B	�x   x   �	�� ��1��� ���	���½�k�b/�&�-�IsY�3����R����¾6�ྺ���	��Z���
Z�	������@����¾�R��1���JsY�3�-�^/��k��½x   x   Nc�˃P��P�fc��U�������`ս@,���4��g�)#������';jW�gy ����o�o����my �fW��';���.#���g���4�;,��`ս�����U��x   x   �\�����\��u2���o�ѻ��&_佹t�y~K�y����������4߾%	��օ� 8���&8�Ѕ�!	���4߾�������{��~~K��t�_�Ż��D�o��u2�x   x   ����ڼ��N��k2��J��Ԫ½�5	�0G:���s��䙾���� ݾ������
�����������
������ ݾ����䙾��s�:G:��5	�ɪ½�J���k2����x   x   ⤼���߼m�%�v���S�½�A��.D��Ԃ����}cоߜ�������!�=S/���7��:���7�<S/���!��������cо����Ԃ��.D��A��½r�����%���߼x   x   ��߼V��p��ܺ��S�E��������޾	5�C���4���F��S�J�Z�O�Z��S���F���4�?�5��޾������I�E����ܺ�ظp��U�Y�߼x   x   �%���p��y��jy
�a�G��J�������8��l.��ZI���`��s���~��:����~��s���`��ZI��l.�9��쾞���J��{�G�my
��y����p��%����x   x   7����ں�Sy
�Y�H�_����ڽ��Q��i���<�o�\��hz�U������]n��\n������	U���hz�h�\���<�i��Q���ڽ�S���P�H�Py
��ں�I���tH��H�x   x   ��½���G�ߎ�� ����M�!�&RG��/m��i���ח�����&?���έ�(?�������ח��i���/m�#RG�D�!����(�㎌� �G�����½�(��7���(��x   x   U@�=�E��K���ܽ�i����	$�'&M�:�w�W���t����1使��ÿ��ÿ1使�r���U���;�w�,&M��	$�]����ܽ��K��;�E�a@�zDҽ0��,���Dҽx   x   �.D��������dU��&�!�e'M���{�E'��Z��.���̿d�տuٿd�տ�̿/��]��C'����{�d'M�'�!�mU����������.D�j��Gs��ٽGs�l��x   x   8ւ�>��V�hl��UG�J�w�5(�����}�ÿ(ֿ�㿜�鿝�鿵�(ֿy�ÿ���8(��G�w��UG�gl�Q�E��<ւ�~�E�����?
��?
������E�x   x   ����#޾���<�O5m���������ÿ�nٿ������,��������nٿ��ÿ�����U5m��<����#޾���
퀾Q�M��0�x&��0�Q�M�
퀾x   x   �hо�9�3s.�]�
n����������*ֿ��tF����������tF���꿹*ֿ�������n��]�3s.��9��hоPg��W����^��mK��mK��^�V���Hg��x   x   ߤ����6cI��rz�4ݗ�����1�̿�"�$���#���b��#���'����"�.�̿����5ݗ��rz�<cI���ڤ����ž�5���q��szx�T
p�wzx��q���5����žx   x   (����4���`�r[���ţ�?뽿�տl��N1����������J1��m���տ?뽿�ţ�q[����`���4�.��:龅���*奾ϕ�uY��uY��ϕ�&奾����9�x   x   ��!�p�F�s�c���zG���ÿ�ٿ������ K�������鿃ٿ�ÿ{G��d���s�p�F���!��� +߾|�¾6԰�f���v��f��>԰�}�¾+߾��x   x   B\/���S�o�~�9w��Lح�H�ÿ��տ'㿱꿫�'㿫�տI�ÿMح�7w��f�~���S�C\/��X�����3ݾ�E˾�M���󼾯��M��}E˾�3ݾ����X�x   x   {�7���Z�RC��(x���I���4�̿H1ֿ�vٿK1ֿ2�̿��I��(x��VC����Z�y�7�����������$�پ%�վ�Ծ(�վ,�پ��⾮�������x   x   �:���Z���~�$����ɣ�-������:�ÿ<�ÿ���+����ɣ�&�����~��Z��:�<!�6[���������|A�`��\��tA� ��������3[�<!�x   x   ��7���S�Qs��_���◿����!!���!�������◿�_��Vs���S���7�(=!����b2��� �7
���b��{���iF ������b��6
���� �b2���&=!�x   x   �`/���F�Z�`� ~z�u��]Ő��1���1��_Ő�u��#~z�W�`���F��`/��!�]�H3���V����h��������h���T���G3�]��!�x   x   d�!�T�4��mI�]��Dm��w�D�{��w��Dm�]��mI�R�4�`�!��]�������y� �/�~��d���������d��0�y� ��������]�x   x   ��8��~.���<��eG�9M��8M��eG���<��~.�7����J�����խ�s���"��.�[e�����p��p����[e�-���v���ۭ����K��x   x   ص���C�f�z�T�!�$�_�!�z�f��C�е��y�7߾M>ݾ��⾣���h���j�����q��)��q�����j��h������O>ݾ7߾|�x   x   �yо�7޾�,��n����������n���,쾻7޾�yо��ž�����¾P˾��پJ����������&r�*r����������J���پP˾�¾������žx   x   �%���1��.���򽾼
����.���1���%���u���B��)�u߰�jX���վ���sJ �'�����Y�����*��vJ �����վhX��v߰�.��B���u��x   x   �䂾ܢ���]��w��������]��Ԣ���䂾O�������X}��ڕ��p��	����Ծn��}����k��f��f��k�r���m����Ծ����p��ڕ�P}������Q���x   x   �GD�H�E���G���H���G�O�E��GD���E���M��*^���x�fc��t���0����վ�I�]i��.�S�,�_i���I��վ+���t���ec����x��*^���M���E�x   x   �T�*���
���
�1*��T����·�= 0��~K�Qp��a��Sn���U��*�پ��������������,�پ�U��Yn���a��Ep��~K�D 0�������x   x   ��½F���\���I�����½
cҽ[���M
���&�{K���x�FՕ� ڰ�lJ˾b��H���� �u��� �K���[��qJ˾�ٰ�AՕ���x�{K���&��M
�\��cҽx   x   c�����p� �p�x���o?��'1����ٽ�I
�50��^��u��c襾��¾�4ݾӤ���0�0����ڤ��4ݾ��¾l襾�u���^�:0��I
��ٽ1��G?��x   x   O�%�zp��%��+H��F���)��̀�|��.�M�����6������(߾)������V�m���V����-���(߾�����6��	���.�M�v��΀��)���F���+H�x   x   h�߼��߼��� H�2���Lҽ���C�E��쀾�e����ž����JS����3!��3!���KS����龌�ž�e���쀾J�E�����Lҽ�1���H����x   x   <�c��}�>�ۧ���Sڽ%k��Y�F ��N��_��I
�� �CB3��6B��K���N��K��6B�DB3�� �I
�\��N��> ��#�Y�2k��Sڽק��c�>�b��x   x   ��hr3�,����ԽV���	`��}����Ǿ����:Z�}Z4��M�{a��p�K�w�M�w��p�{a��M�rZ4�=Z�������Ǿ�}���	`�E����Խ ,��`r3�:��x   x   �>��*��UOӽ���9�d�ަ���zӾQ��S�'��H�:�g�T6������1��@q���1�����P6��D�g��H�I�'�H���zӾ禞�U�d����?Oӽ�*���>���"�x   x   �����Խ؉�3�f�a#��t�۾%E�C24��Z�;�����-��I�����I�1�����4���Z�T24�(E�f�۾W#��)�f�����Խ'����ua��ua�x   x   qPڽ�����d�#$��<v޾K\�	K<�<	h�V ��D�������K��m�ƿ}�ɿo�ƿK������F���[ ��7	h��J<�O\�Kv޾#$����d����`PڽY���J��W���x   x   k�Z`�����ϗ۾*]�^ ?�%5o��y�������r���eп+ݿ����+ݿ�eп�r�������y��(5o�d ?�$]�ȗ۾����W`�k����Z:��Y:�����x   x   ��Y�̀��@Ӿ�G�]M<��6o�鸒��譿�oǿ̑ݿ���a���CF��_������ϑݿ�oǿ�譿븒��6o�YM<��G�?Ӿǀ����Y���������㽓�����x   x   W#��_�Ǿ���64��h�~{���魿~�ʿ���>���4��B��D��5��:�����促�ʿ�魿w{���h��64���c�Ǿ]#��`8U���$���������$�h8U�x   x   �S������
(���Z����4����rǿ1�俢���-��9�k>�7�.������.��|rǿ7��������Z�(������S���r��M�T��30��X$��30�F�T��r��x   x   ��澋`�'�H����B����w���ݿr�����tN�v��w��tN���s����ݿ�w��>������,�H��`���澉��Fe���O[��C��C��O[�Ee�����x   x   $O
�c4�
�g����>���flп»���i��h�i���������glп?�������g�c4�O
���Ӿ�=��d���۠j���_�٠j�`����=����Ӿx   x   �! ��M�&=���	��fS��|3ݿM������-A�Z��Y��+A����R���z3ݿcS���	��#=���M��! �6k��<ž����Z͋�^���a���[͋�����<ž.k��x   x   zL3���a�;�������Yǿ���O�������.Q�������O����]ǿ����<�����a�xL3����0侳��3棾����������6棾����0侌�x   x   =CB��(p�1;���#���ʿt��]���6��w��s��4��d���u���ʿ�#��0;���(p�?CB�T�������־����hҫ�0���1���fҫ������־����U��x   x   <�K�>�w��{���$���
ǿ�7ݿ���0��)���5����7ݿ�
ǿ�$���{��=�w�4�K��'�Χ
��j��;Ѿ��������q����������;Ѿ�j�Ч
��'�x   x   �O���w�=������ X���rпU�ݿ*��*��V�ݿ�rпX������=����w��O��,����,���V⾯�ҾKUʾ)�ƾ&�ƾIUʾ��Ҿ�V�	,������,�x   x   ��K�M-p�ͩ����现�����|ǿ��ʿ�|ǿ���鎰� ��ϩ��Q-p���K��,�\���:�o[�0�߾�&پG־�վG־�&پ6�߾n[�:�a���,�x   x   dHB���a�(B��h��_���߭����������㭨�Y���k��)B����a�gHB�W'����;�Y*���澳�⾞���⾚�ᾯ�����`*�;���Y'�x   x   �S3�{M�>�g�o�����̅��TĒ�ƅ�����q��<�g�{M��S3������
�1���^�J��<.澃.�:{�Cp�A{꾆.�?.�F�澐^�1����
����x   x   V* ��m4���H���Z� h�9Ko�:Ko� h���Z���H��m4�]* �?�����r쾐\�u�߾u���/�p�����p��/�v��s�߾�\⾡r����A�x   x   �X
��k��(�zF4�_<��3?�_<�pF4��(�l��X
�qz��C=��־DѾG�Ҿ�+پi�ᾤ}�"����#��}�f���+پG�ҾDѾ�־B=�uz��x   x   ����	��eV�Qm�Gm�fV������美�ӾPIž���Dǻ�6���G\ʾ�L־��]s�К�Ԛ�Zs뾋��L־F\ʾ8���Fǻ����KIž��Ӿx   x   �e��6�ǾߖӾ��۾��޾ȱ۾ٖӾ1�Ǿ�e������J��i���K�f۫��!���ƾ�վ��k~��q�j~꾝��վ�ƾ�!��d۫�F�n����J�����x   x   y3�����;����9���9��8�������3��񀊾�q��I���#׋�� ��J����x��h�ƾ)L־Z���0��0�\��&L־h�ƾ�x��H���� ��!׋�<����q������x   x   JZ��*`��e���f��e��*`�9Z��PU��T��b[�o�j�i������ҋ��U���Yʾ!*پ��⾭.澗��!*پ�YʾS��ϋ��
���j�����j��b[��T�QU�x   x   �����f��r���������ݒ$��C0�ºC� �_�V���.���֫�&���w�Ҿz�߾~��~��r�߾z�Ҿ)����֫�6��S����_���C��C0�Ւ$�w�x   x   �sڽiսHtӽlսysڽb���������c$��C��j��Ћ�`裾����A;Ѿ#T�+W�k$�,W�)T�<;Ѿ����X裾�Ћ�7�j��C��c$�������U��x   x   ����D��D�������ġ�mP��X�����90�T[�u�����������־�d��#���5��5��#���d��־�������l���T[�:0���?��oP��uġ�x   x   ��>�;�3���>��a��)���G��:��� �$�]�T�]d���:��A7ž�)侤���r�
�J�����G��q�
������)�77ž�:��_d��W�T���$�X����G���)���a�x   x   4��\���"�Z�a����N��\��7U�xp���	����Ӿ�`����̖��'�C�,�F�,��'�ɖ����`��~�Ӿ�	��~p��!7U�N��>��򴡽T�a�&�"�x   x   L�����<Y��{����z.�#q��f����;3&������0�s�E��rV���`�?�d���`��rV�u�E���0�}��$&����;�f��Hq�&z.���{���Y����x   x   ���$M�~����e1��{�l���߾�K�4,�hLJ�\�e�S�|�V���"Ǌ�!Ǌ�W���Y�|�X�e�ZLJ�>,��K���߾]𪾅{�c1���/~��DM����x   x   �Y��|��Z��2�,���>��&,�ܙ�^>�	c������ĝ�&+��Ų��)+���ĝ�����c�K>�ҙ�=,��>��#,����2�(�|��nY��~9�x   x   5w��7���2��|��1ѷ��^����"�L�L�"wx��t������w��������ſ��ſ����w�������t��#wx�`�L���"��^��-ѷ��|��%�2�E��;w��Z�|�>�|�x   x   	�g1�--��-ҷ�������'��V��$������~����ȿzؿ6j�#��7j�zؿ��ȿ�~������$���V���'�����'ҷ�'-��]1�w	�R���1f��W���x   x   {.�f{��A���a����'���Y�)X��ț�������ؿ�q��$��_��`��%���q���ؿ���ț��(X����Y���'��a���A��e{�%{.�%��z�˽~�˽�$��x   x   �q�w����1���"�ߊV�Y���6��>$ƿ�G�����$I��������%I�����G�8$ƿ�6��Y��֊V���"��1�o����q�B�,��_���_�H�,�x   x   #k����߾r��{�L�'��흤��%ƿ����b�?��
��_��a��
��=���b���濊%ƿ㝤�'����L�s����߾'k����f�s�-��x��x�p�-���f�x   x   B�;<Q�U$>�x��������J��c��&�����7$�h�&��7$�����&��c��J㿵����x�D$>�=Q�G�;9����s_��44��,&��44��s_�:���x   x   �1��,��c��z��������ؿ���������&��%,��%,��&����!�������ؿ����}z���c�-,��1��eλ�J����]�CA�CA�ŭ]�I��lλ�x   x   w��WJ����㯤���ȿ�y�L�	��:$�',���.�',�:$����L��y��ȿ䯤�����VJ�l���`侗>���놾n�c�|�U�i�c��놾�>���`�x   x   ��0���e����!�����ؿ�.��á�{����&�$(,�$(,���&�|��ơ��.����ؿ#��������e��0�i�WA;�6��k�r�r�k�7��cA;i�x   x   WF���|�yΝ�e����u�7��~��|��9<$�^�&�;<$�{��z��8���u�d���vΝ���|�UF���E����Xϛ�Չ����Չ�Vϛ����E���x   x   �V�ޑ��H6���ſ<������������������������5��
�ſI6��ᑆ��V�|�(�a��a<վȩ�����*���+������ө��`<վY���(�x   x   '�`��ъ����C�ſ�x�v3�� P����<,����P�r3���x�E�ſ����ъ��`��4�@�2�꾰�žm���(
����d𭾲�ž<��@��4�x   x   w�d��Ҋ�b8���Ŀ�"�ؿ ��{����i��i�}������ؿ�Ŀ�a8���Ҋ���d��9��K�8��ghվ����r���<��	<��y�������^hվ8���K��9�x   x   �`�{���|ҝ�ׅ��!�ȿ!�ؿQV����MV� �ؿ$�ȿՅ��|ҝ�~����`�N�9���C6�R�߾ɾX���h���=���e���W���ɾQ�߾>6���R�9�x   x   ��V���|�Y��@���ڍ�����"2ƿ)2ƿ���ҍ��C���\����|���V��	4��M� 7��<㾋!Ͼ�gþD[���亾�亾D[���gþ�!Ͼ�<�7��M��	4�x   x   FF�u�e���������*$�������C������0$����������w�e�CF�)�(�#� =��>�߾�"Ͼy(ƾ¾	���_e��	���¾{(ƾ�"Ͼ<�߾(=��&�'�(�x   x   ��0�$cJ��c� �x��1���d���d���1���x��c�&cJ���0�!���� ���mվ�ɾjþ¾��¾J�þK�þ��¾¾jþ�ɾ�mվ������!�x   x   ���� ,��3>���L��V���Y��V���L��3>�!,����Lq��Q�7Fվ=�žA�������#^��������þ�ľ��þ����^������F���@�ž8Fվ�Q�Lq�x   x   �F���]�4����"�$�'��'���"�>���]��F���q�O;�������~�����������纾@g��.�þ-�þ<g���纾����
���w����������O;�q�x   x   �;T�tL�l��������]L�V�#�;�޻�0L��)B���؛�$��Z��A�����纾n�����¾u���纾���A��`��$���؛�+B��9L���޻�x   x   �|������X���귾�귾�X������|��]�������h���?���k܉�N������?��᝴�z\��¾¾v\��靴��?����N���l܉�@���^���򋌾e���x   x   54q��@{��?��_����?���@{�4q�W�f�9�_�q�]��c�r���A����������t���zfþ�%ƾ�fþs����������@���	��r��c�~�]�)�_�\�f�x   x   �.��11���2���2��11� �.�,�,�6.�TD4��OA��V��r��׉����𭾔~��u�ȾfϾbϾm�Ⱦ�~��𭾱���׉��r��V��OA�ZD4�7.��,�x   x   �/�=�����9���/�G���n�(��E6&�
JA���c��JΛ�񦱾�žyaվ}�߾h2�}�߾�aվ�ž馱�GΛ�󅾬�c�JA�;6&�.���n��G��x   x   ������ᘜ����*����˽^&���84���]�hꆾ�3�����4վ^�꾿*��s.�v.��*��M��4վ����3��bꆾ��]��84���!&�(�˽5���x   x   %*Y�\�M�k*Y�ʹ|�#v��T�˽�c���-��q_�!|���8���8;q9����#��@�R���@�&����c9��8;�8��|���q_���-��c�_�˽v��̹|�x   x   t�������9�W�|������)���,��f�񏕾Aǻ�V��a���.�(���3�*�9�/�9���3�)�(����a�V�>ǻ������f��,��)������v�|���9�x   x   CS��-�w�r��ϴ���U7?����7���aN����.'��{A���X�t�j���u���y���u�t�j���X�|A��.'���_N�?���+���j7?�����ϴ�ݒr��-�x   x   �-�;�f�������C�C�^���}���0V��i��>�vm_���}�{��7s��������8s��{����}�hm_��>�z�V��h���N���P�C�������{�f��-�x   x   {�r�X���Y�[;F�T5����ƾ4��u�*��S�%�{�L@�������鮿���广����鮿����T@��%�{�xS�p�*�G����ƾT5��J;F�bY�P��V�r���O�x   x   P˴�O���;F��ې�G_̾4�
��R5�d��6��໡�L����ȿ`տ��ۿ��ۿ`տ��ȿG��޻���6��d��R5�!�
�J_̾�ې�<F�Z��J˴����饋�x   x   Z��ғC��6��t`̾.���
;�Uo��+���خ���ȿ�q߿7��/��� ��/��6��q߿��ȿ~خ��+��So�;�7��g`̾�6��ƓC�[��Vý
ի�Výx   x   H9?�˙����ƾ��
�/;�z�r�s闿�M��1�տm��_����k�k����_�m��7�տ�M��o闿w�r�+;���
���ƾ˙��I9?��o���۽��۽�o�x   x   �xü�j��LV5�yo�sꗿ�:����ܿ�T�����a�*��$,"�(���a����T����ܿ�:��zꗿso�HV5�k��nü����:�f��" �c����:�x   x   ����^��Ϛ*��d��.��P��2�ܿ۱ ������h_*�E�/�G�/�h_*������߱ �2�ܿP���.��d�Қ*��^������1y�k�8�������g�8��1y�x   x   �W��#��!S�9;��ݮ�c�տEX������"��0�ؽ8��;�ؽ8��0���"���@X��j�տݮ�5;���!S��#��W��?���l�?�:��*�A�:��l��?��x   x   #��>�X|� ¡�7�ȿ����&���0���;��B��B���;��0�'�������0�ȿ!¡�c|�>���?Qʾ����v�c���B���B���c�����LQʾx   x   �8'��y_��G�����oz߿kc��e��b*�`�8�2B�8E�2B�`�8��b*��e�nc�tz߿~���G���y_��8'��������2�����a��R���a�/����������x   x   ]�A���}���ؙȿ�������/���;��B��B���;��/�������ܙȿ����}�f�A�����x׾Hã�����v?h��?h�����Rã��x׾���x   x   КX����������տ�<����2"�8�/���8���;���8�8�/��2"���<���տ��������͚X���$�����6y��bЗ����v���^З�"y��������$�x   x   a�j�!~��0%����ۿ�	 �����?f*��0��0�>f*������	 ���ۿ4%��%~��f�j��5�TR��׾�G��ԋ��P焾Q焾ڋ���G���׾NR��5�x   x   �v��)����ۿ�?������i�]��(�"�a���i�����?���ۿ���)���v���A���#"�&�������W�����W������"���*"����A�x   x   ��y��*���'���"տ+�g����������g�$�"տ�'���*���y�H�X������G	ξ���W����ݒ��ݒ�d������@	ξ����[���H�x   x   v����3���0�ȿ�߿v��+e��K� �-e��s���߿0�ȿ2������v�W	H��/!������׾�Ǹ�MF������Zj������DF���Ǹ���׾����/!�\	H�x   x   ��j����Y�����q�ȿ��տE�ܿJ�ܿ��տi�ȿ���\��
�����j���A�{��k��h,۾04��X���(��j9��p9��.��W���.4��q,۾i��u����A�x   x   v�X�C�}�@O���ˡ�V访]��II��]��a访�ˡ�7O��J�}�t�X�/�5�������I�׾V5��wꭾ(}���ɟ��b��~ɟ�-}��vꭾP5��H�׾������/�5�x   x   ͒A�-�_�|�FE��4:��m���w���3:��=E��|�2�_�͒A���$��W��)�ξ4˸�/����}��$��Y֟�_֟�"���}��8���4˸�ξ�)��W���$�x   x   �C'�F*>��2S��'d��*o���r��*o��'d��2S�E*>��C'�p�������׾H��!����I��?���ʟ��֟������֟��ʟ�<���I��*���N����׾
���m��x   x   ����1�8�*��h5�� ;�� ;�i5�A�*��1�������ˆ׾'���P����ʴ������<;��jc��w֟�p֟�gc��>;������ɴ�����P��$���Ԇ׾����x   x   �mᾊx��b��g�
����w�
�P���x���m�cʾ��dΣ��ؗ�`����[��Sᒾgl��M:��Xɟ�@��dɟ�I:��al��Tᒾ�[��c����ؗ�`Σ���cʾx   x   ����ڼ���ƾ|̾|̾��ƾ(ڼ�����2P��)
������'���F���넾����ߒ�Ѻ��+��{��{��!��ݺ���ߒ�����넾@��.�������
��:P��x   x   �������lK����cK����������My��6l���c�!b��Ih��v�D鄾gW��3����C��E���F孾O����C��%���qW��D鄾�v� Jh�b��c��6l��My�x   x   sT?��C��[F� \F�ͱC�_T?�@�:���8���:�>�B��R��Ch�b��[���n������������+���+������㚮�r���Y���_���Ch��R�:�B���:���8� �:�x   x   (��ܦ�bp�Ԧ�B���������h�*�}�B���a�e����̗��A������r�;��׾�۾��׾r�;�����A���̗�l�����a���B�e�*��������x   x   t鴽�6��K6��z鴽�qý�۽!+ �]��=�:�F�c�����,���p��ա׾����^w�`w�������ԡ׾*p���������R�c�6�:�]���* �1�۽�qýx   x   կr���f�I�r�踋��嫽.�۽Օ�8�8� l���������l׾I����H�*�,��!!�$��-��H�A����l׾��������l�K�8���?�۽H嫽鸋�x   x   �*-��*-���O�M���^ýFq�M�:��+y�:���Gʾ%������t�$�X�5�ǡA�?�G�G�G�ɡA�U�5�q�$����+����Gʾ:���+y�%�:�Cq�(^ým����O�x   x   �&��??�|����cĽ�y�leN�gR���Y������g\4���P�=�i�O�|�����������Q�|�7�i��P�r\4�ݤ����Y��|R��~eN��y��cĽ'����??�x   x   i8?�z}�hɽ�u���T�NE���̾S,��c)�2N�vLr�+����+���ݠ�饿饿�ݠ��+��)���iLr�2N��c)�B,���̾BE���T�����ɽ��}�?8?�x   x   P���Ƚ�����pW����Pؾ0x�D�9�A�e�����?ܝ�����?��:�ƿ^�ɿ<�ƿ9������Fܝ�����.�e�F�9�Gx�Pؾ����pW����Ƚ�<����c�x   x   p_Ľf���qW�
����޾�3�+�E�5dx�9s��$���+ǿ-ڿ~���������-ڿ ǿ(���Ds��3dx� �E��3��޾����qW�t��b_Ľ��������x   x   �y��T�����Z�޾̋�`�K�"A��DE��4R���ڿN��L�+v	����*v	��L�N��ڿ'R��CE��(A��l�K�ԋ�G�޾�����T��y�ضҽ�#���ҽx   x   hN�+H���Sؾ�5���K��Y���t��@�ǿb�����m����R��T������m���l��E�ǿ�t���Y����K��5��Sؾ-H��hN��y�J��S���y�x   x   V��ϻ̾�{��E��B���u����ʿGZ�b
����&�O�.���1�N�.���&��\
�DZ���ʿ�u���B���E��{�Ż̾V���H�~v���|v��H�x   x   �`��/1�<�9��jx�pH���ǿ�[�]�!5��G/�j;��JA��JA�g;��G/�%5��]��[�ۓǿlH���jx�B�9�+1��`���8��3SC� !�#!�.SC��8��x   x   � �k)�.�e�%x��1W�����:!
�86�O>2�.~A��YK�p�N��YK�/~A�M>2�56�9!
���5W��!x��#�e�k)�� ��O���x�GB��0�GB��x��O��x   x   ���v<N�������#�ڿ���=�PJ/��A���N�[�U�Y�U���N��A�QJ/�?�����ڿ�����|<N�����!ؾ徛�*Zk���F���F�6Zk�⾛��!ؾx   x   Pg4�;Zr�W䝿(ǿ�W�r�y�&�X;��\K���U��{Y���U��\K�V;�x�&��r��W�#ǿP䝿7Zr�Ng4�rS�\J��ܨ����c���Q���c�ڨ��SJ��iS�x   x   ��P�ӝ�����M8ڿ�R���W�.�+PA���N�U�U�W�U���N�+PA�Y�.����R�S8ڿ���֝����P����.F⾕����u���c��c��u������;F⾌��x   x   [�i�S6��L�����`}	�˜���1�~QA��_K�6�N��_K�}QA���1�̜�f}	����D��P6��U�i�(�/�ǜ�z�¾C͖�ޑ{�Fnk�֑{�=͖�h�¾Ɯ�%�/�x   x   f�|��頿�ƿJ�7��՝���.�&;�ބA�ބA�';���.�՝�1��J��ƿ�頿n�|��A�?-�'~ܾ�h���F����x���x��F���h��/~ܾ?-��A�x   x   c�������� ʿ��	�����&�2P/��E2�6P/���&���&	��￪ ʿ����]���ھN�zw�%<�Jj��[�I
�� K}�D
��J�Aj��"<�zw�پN�x   x   ���������ƿG��HV�4w�K��=��=�K�;w�CV�B�翚�ƿ�������$�U�X&�����ʾP#����k��j���[#����ʾ�X&��U�x   x   ������7?ڿ�`�{��W(
��e�\(
�x���`�:?ڿ��������U�_)��:��^Ծ�H����������������v����H���^Ծ�:�d)���U�x   x   �|�=;����� &ǿI�ڿk��Hk�Ik�i��B�ڿ&ǿ���8;���|���N�ZZ&��;�E�׾�/��嚾�X��蘅�񘅾�X��$嚾�/��J�׾�;�TZ&���N�x   x   ��i�$����읿=��gc���ǿ��ʿ�ǿxc��?���읿)�����i���A��{����aԾ�0��"����ˎ�U��S ��U���ˎ�����0���aԾ���{���A�x   x   7�P��hr������U��̃��ڃ��
U�����)���hr�2�P�r�/� 3�D��ʾ�K���暾5̎�E��
	��	��J��5̎��暾�K����ʾD�3�t�/�x   x   �s4��KN���e�o�x�O��2g��O��|�x���e��KN��s4������!�ܾ+q���'��I���Z���U��	���d��	���U��Z��A����'��0q��%�ܾ�����x   x   G��Jz)��9�a�E�-�K� �K�e�E�!�9�7z)�V��6]�U⾋þ�p�����������������E �����y��H ������������������p���þ-U�-]�x   x   8�,?���{G�.���G���8?�(8��4ؾ,Y���	��yՖ��L����x������g����S��V���S��b�������{�����L��zՖ��	��1Y���4ؾx   x   �u��c�̾�oؾ��޾w�޾�oؾs�̾�u��<a���̛�i����}����{�B�x��M}�=��0���U���ǎ��ǎ��U��:��A���M}�I�x�v�{��}��f����̛�Da��x   x   h���\��7ƛ��3ƛ��\��h���G��Ky��lk�O�c��d��rk�9�x�����m����ޚ������ޚ�u�������=�x��rk��d�;�c��lk�Ey��G��x   x   F�N�U;T�>�W�s�W�2;T�0�N��0H�gC��VB�`�F�R���c���{�JC��q혾d���>��($��$$���>��e��u혾JC���{���c�R�\�F�pVB��gC��0H�x   x   ͏���{	������������F!�ڌ0���F�D�c��r��Bǖ�.`���^����ʾ�NԾE�׾�NԾ��ʾ�^�� `��Hǖ��r��5�c���F��0�I!�������x   x   �Ľ�齽j齽�Ľ�ҽ�����?!��GB��Uk�����U�����¾�nܾ�)� ��.��.�%�|)��nܾ��¾@��������Uk��GB�?!�ǩ����V�ҽx   x   �Ǆ��5}�Ȅ��ԗ��4�����dy��QC�W�x�a���,@��8�}���!��i��H&���(��H&��i��!�}��8�:@��N���Y�x��QC�ty���꽏4���ԗ�x   x   �L?��L?�:d�v˗���ҽB{�oH�5���H���ؾ~K�w���/�Y�A���N��kU�
lU���N�Y�A��/�w�K��ؾ�H���4��HH�E{���ҽ�˗��d�x   x   Y4���M����4ѽ�c���Z�����h�Ⱦ�� �����<?��;]���w�����{��n����{��	�����w��;]��<?�~���� ���Ⱦᖾ��Z�`c�&ѽi����M�x   x   ��M�t�����ʽ�=�ƈa��ȟ�p�پû��14��K[�-΀�S<������謹�J���J���謹���R<��(΀��K[��14����R�پ�ȟ��a��=���ʽ������M�x   x   h���9ʽ�Q��^e�oǥ�ln����2�E���t�rӑ�����<���*ʿ��ӿ��ֿ��ӿ�*ʿ =�����gӑ�x�t�=�E����wn�^ǥ��^e��Q�1ʽR���Qt�x   x   �ѽ�=�v_e��䧾b<�6!�F�R�JW��d<���W��U�ӿ<L�����8���6�������>L�F�ӿ�W��t<��BW��5�R�
6!�q<��䧾�_e��=��ѽb���+���x   x   Yc��a�+ɥ��=�ӽ#��iY��Њ�������ʿ?�����������������������?�迈�ʿ�����Њ��iY�׽#��=�ɥ��a�^c��h߽D.Ľ�h߽x   x   ��Z��˟��r�/8!�kY�����<���ԿJ���`��.��?$�ƒ)�Ȓ)��?$�.��`�W���Կ�<�����kY�28!��r��˟���Z�z��������l��x   x   喾��پ���o�R��Ҋ��=����׿� ��Z�e�$���2�rz;���>�pz;���2�f�$��Z�� ���׿�=���Ҋ�c�R������پ喾�&S�`�L�_��&S�x   x   �Ⱦ����E��Z��!�����Կm ����l=*���;��H�H�O�H�O��H���;�r=*����j ���Կ����Z����E����Ⱦ�|��9�L�ֿ'�ٿ'�4�L��|��x   x   �� ��94��t��A���ʿ7���\��>*�E?���O���Z�Q^���Z���O�B?��>*��\�?���ʿ�A���t��94��� �{���K,���bI�=@6��bI�I,�����x   x   j��W[�ڑ��^�����\d�ͫ$�I�;�+�O��g^��f��f��g^�.�O�J�;�ͫ$�Yd����
_��ڑ�W[�f��;������ s�~oK�xoK�) s�����J��x   x   �H?��Հ������ӿ���3���2�=�H���Z�Tf�	�i�Tf���Z�<�H���2��3�����ӿ����Հ��H?��n
��ƾ;Ց�Gtg�F�S�Atg�<Ց�٘ƾ�n
�x   x   !K]��E���G��AX�x��F$��;�8�O��U^��f��f��U^�7�O��;��F$�s�HX��G���E��K]��"�X	�M�������c��c����X���a	��"�x   x   N�w�B����7ʿ;�������)���>���O�՞Z�Fl^�ϞZ���O���>��)����8���z7ʿ=���E�w��d9��3�1Ⱦt�����w��f���w�n���$Ⱦ�3��d9�x   x   �������|�ӿ��������)���;�j�H��O��O�l�H���;��)����������ӿ�������lBL�If�����������o��o���
������Qf�lBL�x   x   A���JY����ֿG���n���I$�]�2���;�5?���;�X�2��I$�v��I�����ֿGY��:���P�Y�t0%�����J��%���c*|���m�[*|�����J�����t0%�T�Y�x   x   �Î�iZ��+�ӿ������8�d�$��F*��F*�b�$��8������1�ӿhZ���Î���`��b-��"�'�ʾ{����;��|Gq�zGq��;������5�ʾ�"��b-���`�x   x   ��� ���<ʿ�_����j�Yd����ad��j����_连<ʿ �����0�`�660��e���Ӿ�3��К��-w���l� -w������3����Ӿ�e�<60�6�`�x   x   n
��x����N��YԿ��进��� �� �������_ԿO��q���q
����Y�;e-��f��׾g�������#�|�Cl� Cl�5�|�����o����׾�f�5e-���Y�x   x   �w�WL��}���i���ʿӗԿ��׿ɗԿ��ʿ�i��l��]L���w�DIL��4%�J%��Ӿ_�������S����l���f���l�M��}���`�����ӾQ%��4%�GIL�x   x   �V]�H݀��㑿EM���Ǫ��L���L���Ǫ�1M���㑿N݀��V]�Sm9�hl��&��!�ʾ�6���������dm���d���d��dm����'����6���ʾ�&��fl�Wm9�x   x   �U?�qg[�ʮt�If���ߊ�����ߊ�Uf��׮t�dg[�~U?���"� ;���RQ���ß�����|���l�Q�d��Bb�M�d���l��|�����ß�VQ����;���"�x   x   m���I4���E��R���Y���Y��R���E��I4����	y
���sȾį��,����>���/w�1Cl�&�f���d���d�;�f�>Cl��/w��>�����į��rȾ���x
�x   x   R� ����*�^K!�}�#�rK!����^� �4��K�ƾ����w���<��A0|��Iq��l��?l���l�,_m���l��?l��l��Iq�G0|�E��u�������O�ƾ^��x   x   ��Ⱦ��پG��^��]�N����پm�Ⱦ½��L����ߑ�����@�w��"o�"�m�{Dq��&w���|�(��6����|��&w��Dq�
�m��"o�(�w������ߑ�-���ƽ��x   x   /����៾.᥾]���2᥾�៾#���}����8���s�=�g�(#c�]f��o�$|��6�����Z����������6��#$|��o�af�.#c��g�/s��8��d���x   x   ��Z���a�L�e���e���a���Z�AS�K�L�6rI��yK�4�S�^c�L�w����]���|����'��˱��ű���'��}���^������9�w�Zc�A�S��yK�rI�u�L�AS�x   x   �z��W�)l�sW�{��� "��'��G6��qK��pg�v����x��T����<���yʾ޻Ӿ2�־�Ӿ�yʾ�<��H����x�������pg��qK��G6��'�&"���x   x    5ѽ��ʽ��ʽ�4ѽN�߽9���Y'���'�0bI���r��Α�v���v�Ǿ?��.	��X�X��W�]�7	��:�ᾂ�Ǿ\����Α�'�r�bI���'�>'�X�����߽x   x   ���5���;��F����?Ľ������ �L�8(��]���4�ƾ<��g)�yY�_!%��Q-��#0��Q-�a!%�pY�h)�J��@�ƾC���>(��/�L�������~?ĽE���x   x   S�M��M�Cit�K����p߽{���#S�0x��g�������e
�w�"�V9�%1L��Y���`���`�y�Y�'1L�#V9�f�"��e
����h���x���#S�����p߽�����it�x   x   �=��2X������ ڽE��ܪc��`�о���1&���F��f����T������f�����T�������f�	�F��1&�����о�ݪc���� ڽ`����2X�x   x   e*X������dӽ����j�nv�����>��c�;��xd��(��DH��XE��M�����������P���ZE��EH���(���xd�t�;�"�����ov��+�j�,���dӽ"���*X�x   x   >}��kcӽc��1o��֬��L𾡈 �8N�$�~�%�������ÿ�ҿ�yܿ�߿�yܿ�ҿ�ÿ�������~�#8N��� ��L�֬�o�G��bcӽ(}�����x   x   ��ٽ&��o�#���x���-(�f�[����f���8ÿ�ܿ��� � ������ ���o�ܿ�8ÿy������O�[��-(��x��6��-o�5����ٽ������x   x   )��u�j��ج�(z����*���b�)���2ӿ9��])���h��v�e���b)�:���1ӿ=�����b���*�z���ج�j�j�1���d轼̽�d�x   x   R�c��y��Q�0(�Q�b���� ���vyݿ�J�?t�!��+��H1��H1��+�!�?t��J��yݿ�������X�b�#0(�Q��y��F�c��� ��c ��c ��� �x   x   5󜾌�⾾� ���[����6����ΐ�����,���:��GD�&�G��GD���:�,���������@��������[��� ����=�D[�ɒ$����ǒ$�O[�x   x   ��о����>N�� ����c|ݿx���W�r�1���D�A\R�؛Y�כY�>\R���D�x�1��W�s��e|ݿ�񱿬 ���>N������оݲ���WS�n�,�r�,��WS�ݲ��x   x   4���;�- �����7ӿ M�
����1�KH���Y��Be�/i��Be���Y�FH���1���#M��7ӿ���/ ���;�=�f���Z����N���:���N��Z��"f��x   x   �:&���d� ���@ÿ3��1x��,�x�D�K�Y�Gi�BSq�@Sq�Gi�O�Y�z�D��,�-x�0��@ÿ ����d��:&��H�^˧�v�x��\O��\O���x�X˧��H�x   x   ��F��0�������ܿ�.��!���:��`R�5Fe��Tq�ru��Tq�2Fe��`R���:��!��.�}�ܿ����0����F�V����̾�.����j�HDV���j��.����̾Q��x   x   �)f�R���ÿ'�V��+��ND�"�Y�4i��Vq��Vq�4i�!�Y��ND��+�Q�'��ÿR��~)f��(��V�=W��W��#�c�-�c�T��HW���V�!�(�x   x   ʻ��Q��e�ҿ�� ����Q1���G���Y�vIe�Li�pIe���Y���G��Q1����� �\�ҿQ��Ļ���9@��d��6̾ҷ���v�%�c��v�̷���6̾�d�y9@�x   x   _�����	�ܿ������R1��QD�BeR�{�Y�~�Y�CeR��QD��R1�������ܿ����_����S��������ﻆ��j��j�����'���������S�x   x   �"������2�߿x������+��:�S�D��H�W�D��:��+���y��,�߿�����"��u�a��<*�$��B)��6|���t�b�d��t�+|��8)�����<*�{�a�x   x   �t��Ȟ��֋ܿ� ���!��,�>2�52��,��!��� �܋ܿȞ���t���8i�(�2����>L˾T��)T��T7e�T7e�4T��]��XL˾���!�2��8i�x   x   t$��H����ҿ�.��3��~�#��Wa�.���~��3��.򿸮ҿI��p$��::i���5�`��ԾY%��ׅ�~ch�Y]�och��օ�C%���Ծe���5�A:i�x   x   .c��yV��l!ÿW�ܿ���T�!�����T����\�ܿo!ÿqV��1c����a���2�K�ڱ׾�y��	����l�{yY��yY��l�����y��ֱ׾G���2���a�x   x   �����X������KÿEӿ#�ݿn��ݿEӿ�Kÿ���Y��������S�xA*�:��>�Ծxz����[sn�XYX�FQ�BYX�Dsn���|z��A�ԾA��{A*���S�x   x   �5f��8��
���������ľ��پ���������
���8���5f��B@�Q�]��0Q˾�'��'����sn�-&X���M���M�K&X��sn�,����'��&Q˾S��O��B@�x   x   G���d�������̐�S ���̐������v�d�G�V�(�#l����/��K��م�l�#YX���M�fJ���M��XX� l��؅�Y���/�����l�K�(�x   x   �H&���;��RN�D�[�7�b�5�b�N�[��RN���;��H&� ���f��A̾ҵ�������V��eh��xY��CQ��M�۷M��CQ��xY�eh��V��瀒�ѵ���A̾�f����x   x   '*�Q��� �$D(���*�7D(�Ǟ �j��1*�n]쾤�̾�b������������t�58e�]��tY�SX��X�SX��tY��]�B8e�	�t����������b����̾�]�x   x   �о� � p��������
p�� ���оy��ڧ��9���%����v�7"j���d��2e�y[h�Rl�.gn�_gn�Ml��[h��2e�a�d�>"j���v��%���9���٧�y��x   x   ���������/���񬾢�����RÑ��g���y���j���c���c��j�݌t��M���΅������ �������΅��M����t�j���c��c���j��y��g��0Ñ�x   x   `�c��k�~Ao��Ao�^k�S�c�n)[�/mS���N��fO��HV���c��v�����4s��������sj��lj��������/s��������v���c��HV��fO�l�N�dmS�S)[�x   x   ��������������I� ���$���,���:�)^O�v�j�������"������:˾�jԾV�׾�jԾ�9˾�����!�����H�j�&^O���:���,� �$�I� �x   x    ڽ1�ӽ�ӽ�ڽf�轀p �����,���N�I�x��'��\L���'̾�������A������F��������澏'̾@L���'��}�x���N���,�����p �ڄ�x   x   ����t��ٓ��}����̽�i �#�$��TS�9V��ç��̾!E�kY�Q��,*� �2��5� �2��,*�A�lY�6E�#�̾�§�GV��US�*�$��i �K̽{���x   x   @X�=@X��������l��� ��
[�
���k]��a;�����(�*@�>�S���a�}!i��!i�z�a�C�S�6*@���(����;�d]��魑��
[��� �m�Q�����x   x   �jB��Y]��Ǘ��޽&�"�h�9 ��x�Ծ"���u)�2�J��j��2������딿GH���딿���}2���j�E�J��u)�#����ԾR ��h���"�޽�Ǘ��Y]�x   x   xQ]��'����׽��"���o��ԩ��{�M��8�?��i��ڈ��R����������6���6����������R���ڈ��i�G�?�.���{��ԩ�3�o���"���׽,(��'Q]�x   x   [�5�׽y+#���s�Qd���C����#��wR����f��č���ƿq�ֿp�� _�r��i�ֿ�ƿč��U�����xR���#��C��0d��z�s�`+#�+�׽E�YÂ�x   x   J{޽��"�� t�����+���H�+�o9`��Ќ�ng��V*ǿN����P�fg�fg��P� ���M�g*ǿ�g���Ќ�T9`�;�+�H�������� t���"�/{޽,���+��x   x   �"���o�5f������ic.��xg�W���;����u׿ޖ���	����E�����E����	������u׿>���n����xg�dc.�����)f���o�"�"���8�Ͻ%��x   x   �"h�bة�@H����+�$zg�E��je�����������p$��`/�,5�,5��`/��p$����#�����\e��7��.zg���+�OH��hة��"h���#���������#�x   x   �������#��=`�L����f�����]<�x�
�/�1�>�N�H��L�L�H�5�>��/�r�]<���忰f��Q����=`��#��������_��e'�J��e'��_�x   x   ��Ծ���~R��Ԍ�ӌ�����G=�<����5��I�
4W�p�^�p�^�	4W��I���5�<��A=����Ќ���Ԍ��~R�����Ծ.\����V�\/�\/���V�.\��x   x   ����?����m���{׿����	�=�5�ߡL�P�^�S�j�!�n�V�j�R�^�ڡL�;�5��	�����{׿m�����ޟ?�����ֿ�ㄈ���Q�}=���Q�℈��ֿ�x   x   y)�$i�y��2ǿ��������/��I���^��n�A�v�@�v��n���^��I���/�������22ǿw�� $i�v)���gu��K1|�\�Q�[�Q�V1|�`u����x   x   �J��∿���MXῐ�	�<v$���>��8W���j� �v��!{� �v���j��8W���>�@v$���	�AX�򖲿�∿!�J��+�"о������l���W���l�����о�+�x   x   q�j��\���ǿ���~ �&h/���H��^�A�n���v���v�E�n��^���H�$h/�z �����ǿ�\��b�j�y�+�&���c�����Red�[ed�����c��&����+�x   x   �<������3�ֿ�X�N��45��&L�x�^��j���n��j�w�^��&L��45�N��X�+�ֿ����~<��ָC�c��D�ξ-�����v��*c���v�&���=�ξ\����C�x   x   ����?��;p�K��+65�P�H�M=W�K�^�M�^�N=W�P�H�)65�E��<p�G��񒵿���ܟW�u��� �Yq��6S���%h��%h�;S��`q��� 龈��ڟW�x   x   ����F���p�q� P��k/���>�� I���L�� I���>��k/�(P�q��p�F������g�e��,������ཾ����7eq��4a�5eq������ཾ�����,�o�e�x   x   �V��JG����[�^$��{$���/��5���5���/��{$�Z$�[�"��JG���V��Utm��q5�!2���˾���k|�{�_�|�_��k|�����˾#2��q5�Qtm�x   x   ����p�����ֿ�����	�w����خ���s����	������ֿq��������um��e8����K*վ�����P��Һa�I�U�ĺa��P������?*վ����e8��um�x   x   E��(���?ǿQbῼ���s��$F�F�p������Tb�Bǿ���H���e�Gt5����Zؾ1��䆾�d�x�P���P��d�䆾 1���Zؾ��@t5���e�x   x   �A���c��?����=ǿg�׿���忱�y�׿�=ǿ0����c���A���W���,��4��,վ�1��z,���`f�r�N�9KG�a�N��`f�f,���1���,վ�4���,��W�x   x   ��j��ꈿ���[y������v���v�����Dy������ꈿ�j��C�ۉ����� ̾k���冾,af�gXN��
C��
C��XN�Jaf�冾k���� ̾���؉��C�x   x   ��J�X5i�:&������1Ó�;"��Ó�����@&��E5i���J���+����+龎罾����R���d���N��	C�O?��	C���N��d��R������罾+�����+�x   x   C�)��?�*�R��T`���g���g��T`��R��?�[�)�w6�J6��ώξy��jő�vp|��a�$�P�uHG��C��C��HG�5�P��a�rp|�Vő�y��юξf6��r6�x   x   �������#���+�`y.��+�k�#������%��=оeo������W���iq���_�T�U�8�P���N�WQN�r�N�2�P�5�U���_��iq� X�����Qo��3оZ��x   x   �վ{���g��/��������g����羞վ�鿾_��������B�v��(h�k3a���_��a��td��Sf��Sf��td���a���_�=3a��(h�-�v�#�����9����鿾x   x   ���奄����Ͳ�����奄���l��	����D|�O�l��kd�h+c�^!h�\q�n^|�<H��چ��!��چ�9H��Y^|� \q�k!h�l+c��kd�	�l��D|�����l��x   x   KCh�s�o��'t��'t�+�o�@Ch�.1_���V���Q�D�Q���W�]cd��v�nL��.������z磾?!��8!���磾���#���rL��ͫv�Wcd�޵W�=�Q�K�Q�$�V�1_�x   x   ��"�#�G#�#�-�"���#�fw'��h/�}"=���Q���l����������d���н���˾�վzCؾ�վ��˾�н��d����������X�l��Q��"=��h/�ow'���#�x   x   1�޽�ؽ�ؽ!�޽$���0S�s`/�[�Q��)|�z���TX���sξ�龭���S$�������X$�»���龤sξ7X�������)|��Q�m`/�S������x   x   ٗ��=��[ٗ��A���нٿ�:h'���V� ����l�� �Ͼ�����Tu�z�,�#_5�xQ8�$_5�~�,�@u����!����Ͼ�l��4���2�V�Eh'����н�A��x   x   �g]��g]�Ђ�\7���코�#��_�*W���Ϳ�J���!���+���C��W���e��\m��\m���e��W��C���+��!�o��Ϳ�W���_���#�r�콜7��$Ђ�x   x   ~)B�f]������A޽��"���g�֟��Ծ���I)���J�uXj�4���㍿�Ĕ�� ���Ĕ��㍿*��qXj�͝J��H)���O�Ծ֟���g�;�"��A޽a���_]�x   x    
]������׽��"��qo������<���b?���h������(��-l���T���������T��.l���(��������h��b?����e<羭���ro���"��׽����	]�x   x   ,�����׽0�"�m�s��3������Z�#��=R��J䚿�]����ƿ��ֿӭ�z!�խ࿪�ֿ��ƿ�]��:䚿���=R�{�#������3��O�s��"���׽���z���x   x   V=޽��"�[�s������V��s}+�\�_�B���)9����ƿ)�����-�HB�GB�-�����Ί�ƿ<9��1���@�_�f}+��V�����n�s���"�:=޽j���)���x   x   t�"�ato��5��WX���2.��8g�늓�X���;׿�S���	������ג������%�	��S���;׿X������8g��2.�>X��|5��Vto��"���0�Ͻ4��x   x   O�g�(���>���+�:g�?ꕿ�2��������W��A$��-/���4���4��-/��A$��W�����Ῥ2��1ꕿ:g��+�M��.���A�g��#������#�x   x   �ڟ�iC羏�#���_������3���U��A���/�I�>��{H���K��{H�L�>��/�:����U��3��匓���_���#�^C羜ڟ���^��>'�(��>'���^�x   x   ��Ծ}���DR������[�������x���5���H���V��a^��a^���V���H���5�x�����῟[�������DR�z����Ծc7��`�V��7/��7/�`�V�c7��x   x   ����k?�!����>��sA׿���g��خ5��cL�b�^��Qj�Tn��Qj�d�^��cL�֮5�m�����iA׿�>��$����k?���� ����f��G�Q���<�D�Q��f��$���x   x   �R)���h�\뚿Q�ƿ�[���[���/���H��^��ln��v��v��ln��^���H���/��[��[��d�ƿZ뚿��h��R)�v]�:P���|��gQ��gQ��|�3P���]�x   x   ��J�轈��f��fΊ�	�HG$���>���V��Tj���v���z���v��Tj���V���>�LG$���	�Z��f�����J�q��Ͼ䖾^�l�ǛW�W�l�䖾�Ͼm�x   x   �hj��2���ƿ�������+5/�ڂH�h^�6Yn�h�v�i�v�:Yn�h^�؂H�)5/���������ƿ�2���hj���+�����TF������Yd�Yd�����^F������
�+�x   x   .�� x��p�ֿ�4�"���4���K��i^�8Xj��qn�4Xj��i^���K���4�"��4�i�ֿx��'����C��v�/bξ}���v��/c��v�}��(bξ�v�x�C�x   x   c�b�����K�t��5���H�#�V�Z�^�\�^�$�V���H�5�n��K���࿈b��k�jW�Oa��辺d��fV���;h��;h�lV���d����aa��jW�x   x   Ҕ����2��K�$��8/��>���H�WlL���H��>��8/�%$��K��2���Ҕ�˻e�.�,�4����Խ�ȑ�ڊq�Dba�؊q��Ǒ��Խ����.�,�ӻe�x   x   /��I��z��87�����L$�˧/���5���5�Ƨ/��L$����27����J�� /���9m�)K5�:���˾�&���|��`��`��|��&����˾<�"K5��9m�x   x   Ԕ�f��ֿ߰������	��b�����������b���	�����ֿ߰f���Ӕ�;m�b>8�{�Sվ����o��b��.V�b��o�����Hվ�{�d>8��;m�x   x   $󍿥}����ƿg%�{h��m��� �� �i��yh��k%῿�ƿ�}��'�e�e��M5�l|��Nؾ/?��,��_�d��JQ��JQ�d�d�C��<?���Nؾj|��M5�_�e�x   x   Z��:��p���ǿ3O׿���{g忦��EO׿�ǿ�o��:��]���qW���,���� վ@���O��|�f�5RO�b�G�#RO�`�f��O��@��� վ����,��qW�x   x   auj�ƈ�{���K���i���C���C���i���J������ƈ�Wuj���C��g�������˾Q��8����f�)�N�D�C�@�C�M�N��f�;��Q����˾r����g�ƑC�x   x   `�J��h����#�������2�������4��������h�W�J�l�+�W~�w�E۽�w*���q��s�d��QO�m�C���?�g�C��QO�z�d��q���*��P۽�~�R~�`�+�x   x   _`)��|?�YR��`�qSg�sSg��`��XR��|?�w`)�K����mξjl���̑���|�2b�5IQ���G� �C��C���G�FIQ�9b���|��̑�il���mξ#��F�x   x   ���B���#��+��H.�+�+���#�]��ĩ��r�3�ϾR������*[��D�q��`��+V�LEQ�`KO�"�N�>KO�GEQ��+V��`�\�q�3[�������Q��(�Ͼ�r�x   x   n�Ծ,_��#���z���z���#��L_�9�Ծf���/_��K�����v��>h��`a�`�/b��d�t�f���f��d�Db�)`��`a��>h���v�`���	_��^���x   x   �f���O��/���O��i����H���s��'|�
�l��_d�t0c�V7h���q���|�g��G����D��2���g����|�Ёq�c7h�z0c��_d�þl�j|��s���G��x   x   �h�@�o���s���s���o��h�s�^�T�V�9�Q��qQ���W� Wd�C�v��O��q������i���e/��^/���������f����O��)�v�Wd��W��qQ��Q���V�P�^�x   x   0�"�5�"�0#�$�"���"���#�P'� D/�� =�iQ�W�l�����s��$X���Ľ���˾�վ�7ؾ�վ��˾�Ľ�X���s��8����l�iQ�� =��C/�'P'���#�x   x   4a޽��׽��׽$a޽/��.��/1��;/��Q�?�{��ܖ��:���Rξ<�����r�Ll�Dl�w�2���8�辗Rξ�:���ܖ�v�{���Q��;/�1�?�����x   x   諗����(���N����Ͻj���@'�i�V��a���G�� �Ͼ����'k�4S���,�{85�2*8�|85���,� S�(k�������ϾuG��
b����V�A'�u����ϽM��x   x   � ]�J ]�$��������ԟ#��^�b2��$����O����b�+��xC��WW�V�e�,"m�6"m�H�e��WW��xC�J�+�����O����=2����^��#�������B���x   x   :�<��`W����MKٽ�)���b�s���2о����%��QF��ee��M���犿���L�����犿�M���ee��QF���%���3о�s����b�D)�?Kٽ�����`W�x   x   �XW�hu��ԯҽs5��4j�量�%⾉D�,;�:�c�Ҽ��3Η�����8l����������:l������4Η�м��F�c�",;�mD�r%�量!5j��5��ҽ�u��zXW�x   x   ������ҽrZ�Un��G����7 �V�M��$~�M}���x��=q¿�ѿV�ۿ�%߿X�ۿ��ѿEq¿�x��>}���$~�g�M�T �'���G���Tn�WZ�w�ҽ������~�x   x   Gٽ�5��Un�ƃ�����\�'���Z�X���{��v�¿@$ܿ-U�F ��A��A��F �-U�0$ܿ��¿({��K�����Z�M�'�����ڃ��Vn��5��Fٽ8�����x   x   e)�g7j��I��j���F*�3b�
F��]����ҿB��Ϲ�b��<����:��b��Թ�C��k�ҿ]��F��<b�F*�Q����I��[7j�n)�߬��c˽���x   x   �b�h�z�ﾈ�'��b�����y����ܿ�� ����pw ��+�3�0�6�0��+�kw ������ ���ܿm�������b���'����m��b�KJ �V �[ �>J �x   x   �w��=,�P ��Z��G�����+Q���!I�@}+��:��C�}�F��C��:�A}+�I���+Q࿸���G���Z�Q �2,��w��=lZ�� $��w�� $�FlZ�x   x   �:оJ��M������`����ܿ�����_1�`�C��Q���X���X��Q�^�C�_1��������ܿ�`�������M�J��:о�G��@�R�vX,�zX,�=�R��G��x   x   U��|4;��.~������ҿ� �8K�D`1��^G�Y�'ld�uTh�+ld�Y��^G�B`1�;K�!� ��ҿ�����.~�z4;�^��ܻ�����\N��Y:��\N����ܻ�x   x   �%��c�5����¿5����ր+�1�C��Y�`lh�-qp�+qp�^lh��Y�2�C�Ԁ+����2��"�¿5�����c��%����y`��~x��O��O�~x�r`��ě�x   x   9^F��ą�݁��@.ܿ(���| �0:���Q�tod��rp���t��rp�qod���Q�2:��| �,��6.ܿЁ���ą�@^F�[$��H̾^放�j��
V��j�`放�H̾V$�x   x   ue��ח�x|¿�a�-���+��C���X�rYh��tp��tp�vYh���X��C��+�(���a�|¿�ח�tue��`(���D��������c���c�}���N������`(�x   x   gW��d˦�o�ѿN �j��˵0� �F�P�X��rd�Oqh��rd�P�X��F�̵0�p��N �f�ѿ]˦�bW��t�?����˾����v���c��v� �����˾�c�?�x   x    󊿶y����ۿ|J�n����0�ɟC��Q��Y��Y��Q�ʟC���0�g��|J���ۿ�y���o,S�O��71�ď��d̆��mj��mj�j̆�͏��C1�]��n,S�x   x   ٰ���
���6߿RK�c��+�P$:��C�cgG��C�M$:�+�l��SK��6߿�
��Ұ��J6a�M�)�������������u���e��u��������{���M�)�P6a�x   x   F������ۿ�P ���6� �ȇ+��h1��h1�Ň+�?� ����P ���ۿ��L��A�h��>2�ԅ�1˾KC��Ϩ��f�f�ڨ��VC��$1˾օ�z>2�<�h�x   x   ����$}���ҿci�_��h�HS����SS�d�^��ii�ҿ%}������ΐh�R%5��
�/eԾ�T���;��+mi�]%^�mi��;���T��&eԾ�
�V%5�Րh�x   x   �����Ц���¿8ܿ���� �J�F��� ����8ܿ��¿�Ц������:a��@2���
���׾欩�	��REm���Z���Z�^Em���񬩾��׾��
��@2��:a�x   x   y\���ޗ�늮�i�¿��ҿ3�ܿ�b�*�ܿ��ҿk�¿ۊ���ޗ�|\���3S���)�z���gԾӭ���}���o���Y�s�R���Y��o��}��׭���gԾ�����)��3S�x   x   Ɓe��̅��������n��1)��F)��zn������.����̅���e�z�?����ͯ���5˾uW��*����o���Y�)dO�.dO���Y���o�/��qW���5˾ï������?�x   x   �kF���c�C~�暉��U��U���yU������C~���c��kF�k(�{��;�w��HG���=���Fm���Y�}cO��L�wcO�i�Y��Fm��=��UG�����;�v��j(�x   x   k�%�AE;��M��[��%b��%b��[�ڧM�,E;���%��.�����˾z���a���T����ni���Z�1�R�laO�baO�P�R���Z��ni�T���Q���y����˾���.�x   x   >���Y�g �}�'�y[*���'�K ��Y�H��\��eX̾�������Qц��u�f�4#^�)�Z���Y�,�Y���Y�"�Z�#^�f��u�[ц�󞘾���bX̾���x   x   bRоfG�]���������e�ﾁG�4Rо�0o��;������v�Kqj�ыe�pf�Nei�;m��o�D�o�;m�]ei�~f���e�Qqj���v���D�o���x   x   ��	���b��V����b��%	������^X�����.�x�ޕj�p�c�d�c�jj��u������3�����Vs������3�������u� jj�k�c�t�c���j�l�x����?X��x   x   c�p[j�C|n�v|n�3[j��c�V�Z���R��lN��O�CV�7�c�"�v�4Ɔ�����8��OG��띩�䝩�`G��8������7Ɔ�	�v�2�c�eV��O�blN��R�6�Z�x   x   �A�XP��u�FP��A��_ �(2$��d,��`:�'O���j�)���h���䃫�����˾�PԾO�׾�PԾ�˾����ك��l���?���|�j�$O�a:��d,�02$��_ �x   x   ;jٽ+�ҽ�ҽ0jٽh��= �����\,��[N��vx�Xߔ�w�����˾@澀����x�l�
�d�
��x�����;���˾[���_ߔ�0wx��[N��\,����M ����x   x   ���抍�$���-��v˽� �]#$���R�Q���5X���;̾��������E�)�o,2��5�n,2�H�)��������� <̾X��^�����R�g#$�� �uu˽�-��x   x   �nW��nW���~�_#��ٴ�%K ��hZ�+C��rӻ�p�����T(��?�7S�o!a�*xh�6xh�e!a�<S�1�?�T(������kӻ�
C���hZ�3K �2�罚#���~�x   x   �&3�ܡL�3/��W�Ͻ��M�Y�a���Ǿ�; �����E>�y\��Cv��P���ȋ� ��ȋ��P���Cv�}\��E>�����; �%�Ǿv��Y�Y�И�G�Ͻ�.��֡L�x   x   ��L��Ά�7`ɽl��X`���W�ؾ~���=3��$Z��!���y���П�P��Pa��Na��T���П��y���!���$Z� >3�g��9�ؾ��Y`�#l�[`ɽ�Ά���L�x   x   �)���^ɽ�}�r$d��㤾�0����D�~Bs�8��+���@���ɿ��ҿ
�տ��ҿ�ɿ�@��1��.��mBs���D�.��0��㤾V$d��}��^ɽ�)����r�x   x   �Ͻl�F%d����a��bU ��yQ������a��IY����ҿ4�z���X*��V*�����6���ҿTY���a��젃��yQ�PU �p�����`%d�l�	�Ͻ�ɠ��ɠ�x   x   Ø�8[`��夾����"�;X�w��yͩ��ɿ��翉� �;���������;��� ����ߕɿzͩ����(;X��"���뾂夾,[`�ɘ�GF޽�0ý^F޽x   x   g�Y������4�sW ��<X�K���K���dӿN���
��pS��R#�t�(�v�(��R#�jS���[����dӿ�K��K���<X�vW ��4�����_�Y�/�gz��pz��#�x   x   w"����ؾ���}Q�L��!M����ֿ������f�#�
x1�F`:�[v=�D`:�x1�g�#���������ֿ*M��O���}Q�����ؾ"��!)R��`�����`�,)R�x   x   ��Ǿ����D�n����Щ�lgӿǸ�����
E)�޶:�^�G�<RN�<RN�[�G�ܶ:�E)����ø��igӿ�Щ�r�����D������Ǿ�Ջ��K�$ '�( '�	�K��Ջ�x   x   �A ��E3�Ls��f��>�ɿ4������7F)��=�2�N�gAY��\�jAY�4�N��=�4F)����<���=�ɿ�f��Ls��E3��A �CԴ������H��5���H����EԴ�x   x   ����/Z�����`��<��Š�ǽ#���:���N�O	]��d��d�M	]���N���:�ǽ#� �6�翜`������/Z�����������Cr���J���J��Cr�������x   x   �Q>�9)���"��m�ҿ�� ��X� }1���G��DY���d���h���d��DY���G� }1��X��� �d�ҿ�"��:)���Q>�?�	���ž�l���g�T�S��g��l����ž8�	�x   x   �.\�򂑿�K��(翍A�6Y#��f:�!XN���\�)�d�,�d���\� XN��f:�3Y#��A�/翧K�������.\�"�?"뾇 ��݂��c�c�ۂ��� ��I"�#"�x   x   Vv�ܟ�a'ɿĢ�������(�Y~=��YN��GY��]��GY��YN�X~=���(��������X'ɿܟ��Uv���8�e����Ǿ�^���	x��]f��	x��^����Ǿ`����8�x   x   �[��/��b�ҿ�:���%���(�^i:�ʑG�z�N�|�N�̑G�`i:���(��%��:��i�ҿ4���[���RK�����m�B���:C���o��o�AC��N����m�����RK�x   x   �ԋ��o��V�տL<��n��r\#�ҁ1��:���=��:�́1�o\#�v��N<��Q�տ�o���ԋ��X��$������5��6Ӕ�+,}�8�n�$,}�(Ӕ��5�������$�
�X�x   x   i���p���ҿr��� E��]�R�#�6N)�/N)�P�#��]�E�k����ҿ�p��o��<�_��,�@��Hyʾ���'ᅾG�r�E�r�5ᅾ��UyʾB���,�6�_�x   x   �֋�{��u,ɿ~#翕� ���*��f��2������ ��#�u,ɿ|���֋���_���/�+�|�Ӿ)��� \���y���n��y��[�����u�Ӿ-���/���_�x   x   _��C៿�R����ҿ�翃���6���3����������ҿ�R��<៿	_��`�X�>�,��]�־�0���͐�r�~���n���n���~��͐��0��]�־�8�,�^�X�x   x   �_v�����{+��lk��%�ɿpvӿ��ֿfvӿ8�ɿmk��k+�������_v��YK�v�$����"�Ӿ�1��ab��(;��*�o�I�i��o�#;��Sb���1��'�Ӿ���x�$��YK�x   x   e:\��0��W��Pr��-ީ�\��\��(ީ�<r��d���0��^:\�R�8��������E~ʾ򠨾�ΐ��;��:p�ָg��g�Mp��;���ΐ�젨�<~ʾ�������U�8�x   x   �^>�@Z��_s�௃�J ��'Y��B ��쯃��_s�@Z��^>��""�����w�P<��- ��X^����~���o�{�g�Qe�w�g�q�o���~�S^��: ��U<���wᾛ���""�x   x   ���U3���D�x�Q�TTX�KTX�}�Q���D��U3���~�	��1�͏Ǿ���Hؔ�䅾�y��n���i�ٶg�Ƕg��i���n��y�䅾;ؔ����ˏǾ�1�t�	�x   x   RN ���E.��j ���"��j �,.���]N ������ž�+���f��~H��02}���r��n���n�g�o��p�i�o���n���n���r�72}��H���f���+����ž���x   x   ��Ǿ��ؾ.R�����3R徱�ؾ��Ǿu派>��?w��h���0x���o��n���r�y�6�~�6��)6��$�~�&y���r���n��o�x�y���Aw����x派x   x   �5���
��q���c��u����
��s5��w勾����sVr��g��c�O`f�J�o�$&}�C܅�HU���Ő�WY���Ő�QU��6܅�3&}�Q�o�U`f��c�qg��Vr�����_勾x   x   %�Y��}`��Id�!Jd��}`��Y�CCR��K�C�H���J�]�S��c�[x�&>���˔�(��?���M#��G#��D���)���˔�'>��Gx��c�m�S���J��H�9�K�)CR�x   x   &��ƅ������_���(�tq�g,'�M�5���J�V
g�b~��W��ł���'���hʾ��Ӿ��־ȭӾ�hʾ(������W��t~��8
g���J�e�5�h,'�|q��(�x   x   �н,�ɽ��ɽ�н�d޽��������$'�W�H��=r�Tf������vǾU\ᾀp��
���������p��O\�wǾ���Vf���=r�.�H��$'��������e޽x   x   ]?��lㆽ�?���ޠ�vBý���Wc��K����s����žN������$��,�Tz/��,��$�����\��žY�������K�`c������Aý�ޠ�x   x   @�L��L���r��Ԡ�4N޽9�&R�Jы�B̴�V��~�	��"�;|8��AK�Z�X�m�_�y�_�U�X��AK�H|8��"�|�	�q��C̴�/ы��%R�A�wN޽�Ԡ�3�r�x   x   Y%�$�=�B�����½as�^�L��W��5���h����3��BO���g�!{������������!{���g��BO��3����h�J���W��p�L�=s���½� �=�x   x   ��=���z��P������R��-��8˾)1��&(�d�L���p�𖈿���/���b���`���2���������p�r�L��&(�1��7˾�-��%�R�����P���z�q�=�x   x   ���BO��q���U�������־�a��98�g�c�F������� ��������pſ:uȿ�pſ{����������A���T�c��98��a���־�����U�P��:O��	����b�x   x   ��½�����U��i����ܾ��?D�,�v�'R�����טſ̌ؿ�濲)�)���Όؿ͘ſ!���1R��+�v�4D�|���ܾ�i����U������½����њ��x   x   �r� �R�F����ܾ'_�uXJ��C��P��P弿��ؿ�x�mM��h���
��h�mM��x��ؿC弿P��D���XJ�/_���ܾ;����R��r��@ѽ�޷��@ѽx   x   ��L��0��Z�־w��YJ��X��q5���ƿ��f���O��}��S��S��}��O�g�����ƿl5��{X���YJ�w�m�־�0����L�$���h齱h���x   x   s[���=˾je�D��E���6��7>ɿЉ��	�@���l%���-�?W0��-��l%�B���	�͉�9>ɿ�6���E��D�ke��=˾{[��	�F�K�����H���F�x   x   ���5��?8���v�w���ƿd��I�8����-�?�9�ҩ?�ҩ?�=�9���-�<��I�b�ƿs����v��?8��5����e���GB�VF �ZF ��GB��e��x   x   s��-(�@�c�	W��C꼿.��	�L���0���?�o�I�n�L�q�I���?��0�I���	�6�G꼿W��4�c��-(��s�^@��'�w�(~A���/�*~A��w�`@��x   x   ����L�h���魮�� ٿک�Z��>�-�&�?��M��T��T��M�(�?�?�-�\��ة�� ٿﭮ�m�����L���a�־4���P�j�.LF�%LF�]�j�1���p�־x   x   �)3�F�p�����¡ſ��oT�|q%�"�9�E�I�>T���W�>T�D�I�!�9�zq%�rT��񿾡ſ����A�p��)3�Ņ��]��e6���c�^�Q���c�d6���]�����x   x   �PO���������ؿcS�����-�-�?���L��T��T���L�-�?��-���^S���ؿ��������PO�A���0�>���=]���(d��(d�;]��I����0�D��x   x   ��g����u���%&��o�=[��^0�|�?��I��M��I�{�?��^0�>[��o�"&�m��������g�<�.�>��t¾Ɩ�6|�(l�/|�Ɩ�t¾=��:�.�x   x   �4{�&��~ſ�8��
�D\�;�-��9�j�?�j�?��9�?�-�D\���
��8�~ſ*��4{���@��|���۾)q�����b/z�e/z����8q����۾�|� �@�x   x   =����Ť�k�ȿ`:�q����u%��-�D�0��-��u%����q�b:�g�ȿ�Ť�6���9~M������>��̆���腾�9��腾����6�������8~M�x   x   Nͅ��Ƥ��ſ*濲V�Y�Y��������Y��Y��V�{*��ſ�Ƥ�Tͅ�F5T���%�� ��˾�ԥ�����F���F������ԥ��˾� ���%�@5T�x   x   ����>ş�:���ʞؿB�񿵯��	�0Q��	����C��͞ؿ9���@ş�𶃿�6T��D(����܂Ծ`���疾����JP�������疾^��قԾ����D(��6T�x   x   �;{��$��������ſ�ٿ�(翮��(��ٿ��ſ�����$���;{�X�M���%�����׾M���:������t���t������:��N���׾����%�V�M�x   x   �h�ʥ���������c����"ƿ�Mɿ�"ƿs����������ϥ���h�u�@�V��y� ���ԾZ�����S����Y��,���Y��T������W����Ծ� �X��v�@�x   x   �[O���p�a���a������D���D������a��k����p��[O�{�.�ʂ�v���˾d��`<����������B���B���������j<��`���˾n��ɂ�}�.�x   x   �53���L��d�1�v��Q���e���Q��?�v��d���L��53����/���۾&���}٥��ꖾ	��SZ���B��x����B��PZ��	���ꖾ�٥�,�����۾-����x   x   ?��=(��Q8�G)D�pJ�pJ�J)D��Q8��<(�N��{���?�%¾%y��Z���*
�������u��4��dB��[B��6���u����+
��M���%y��"¾�?�r��x   x   Ί��C��u�O �dr�b ��u��C���9�־�l��t���XΖ�캋��셾�H��Q��Bt��`X����jX��>t��Q���H���셾򺋾YΖ�j����l��X�־x   x   (��V˾�־��ܾ��ܾ	�־$V˾�'���Q������@��e��%|�-6z��<��F��'�����������������0����F���<�36z��$|�e���@������Q��x   x   am���D������b��������D��Tm���t��N�w��j���c��1d��,l�80z�S煾b���▾�4��T���4���▾T��[煾<0z��,l��1d�q�c��j�K�w�xt��x   x   �M�^�R�/�U�d�U�;�R��M���F�\B���A��VF���Q��*d��|����� ���?ͥ����)���%������@ͥ�#��������|��*d���Q��VF���A�1\B���F�x   x   ������ �=�����f��~R ���/�~OF���c�Z��L����h��t��% ˾�rԾj�׾�rԾ ˾t���h��R���Z����c��OF���/��R �s�����x   x   �ý�p��bp���ý�]ѽ�齒���K ��~A��j�j1��2z���h¾��۾6��8� �������=� �0���۾�h¾z��j1��(�j��~A��K �u����(^ѽx   x   x����{�����ڮ���﷽u�>���FB���w����S���"����q������%�`4(���%�����q����"��S���򚾥�w��FB�M��0u�D﷽ۮ��x   x   ͕=���=��$b������Hѽ{����F��a��X9��l�־�}���=�.�l�@�GlM�X!T�c!T�FlM�l�@�A�.����}�|�־[9���a����F�|���Hѽ����2%b�x   x   �|�+��p�m���f�,�=��Ђ��
���d߾�o
��%�E�?�i�V�Ȍh�/�s�9�w�,�s�ǌh�i�V�N�?� �%��o
��d߾��т�@�=��f�b��=p�+�x   x   �+��(d�`��=Q���A��R��-��3�� ��S<�;a]���{�Q6��`��q���p���b��T6���{�-a]�+S<��� �����R����A�NQ�;`���(d��+�x   x   �p��^�����ZD��ٍ���ľI�6�(�FQ���y�����q��8D���_���%���_��4D���q�������y�2Q�1�(�[���ľ�ٍ�}ZD����^���p�_�M�x   x   ��Q�[D�ax���cʾ j	���3���a����8-���B��#�ƿ�ӿ;yٿ8yٿ�ӿ&�ƿ�B��6-�������a���3�j	��cʾex��<[D�Q����R���R��x   x   �e��A��ڍ��dʾ�{�39�:�l�!���i&���ƿ�FݿK��˶��B���̶��J�Fݿ�ƿe&�� ���7�l�39��{��dʾ�ڍ��A��e�����b�����x   x   �=��T���ľ�k	�A49��p�m�������ӿ�>￫�L�D��E��L����>￣�ӿ���m���p�>49��k	��ľ�T��	�=��Y��ڽ�ڽ�Y�x   x   �ӂ���s���3�U�l�n���j����ڿ����%�������A} ������'��������ڿ�j��n��P�l��3�t�����ӂ��w9���`������w9�x   x   ������}�(���a� �������ڿ�����+��L���(��-�
�-���(��L��+������ڿu���������a���(��������Yw�.�7�����*�7��Yw�x   x   �m߾w��8Q�w䈿�*����ӿ9����,��� �..�Y�6�R�9�Y�6�..��� ��,�4�����ӿ�*��r䈿'Q�y���m߾�����j���9��!*���9���j����x   x   |v
�G\<��y�g3��t�ƿE���O�C/.��9�3�?�3�?��9�C/.�O���E�m�ƿh3���y�S\<�vv
���Ⱦ{/����b���B��B���b�y/����Ⱦx   x   ��%�km]�\珿�J��BOݿ�����i�(���6���?��
C���?���6�h�(������FOݿ�J��Z珿am]���%��$������E��,�a��-R�'�a��E��y���$��x   x   u�?�U�{��z��A�ƿ�Q�;��.��9���?���?��9��.�=��Q���E�ƿ�z��W�{��?�{���\־Z`�������h���h����d`��]־x��x   x   h�V��?��O���ӿ����ܣ��� ��.�H�6���9�H�6��.��� �ޣ������ӿO���?��e�V���#�����7��F��𙂾=nw�홂�B��$��������#�x   x   w�h�*%��-l���ٿ���Ǥ�D
���(��3.��3.���(�I
�Ǥ�����ٿ1l��.%��z�h�J4��
��A׾	���XV����^V������A׾�
�J4�x   x   B�s��Ɨ�W3��\�ٿ����.T����1T�� �5T����,T�����^�ٿU3���Ɨ�6�s�(P@�O�>���c������,����}��)��������c��E��O�$P@�x   x   4�w�{Ǘ�{n���ӿ���J��r3�n3�J���
�ӿ|n��zǗ�@�w�$�F����
N���ξtɯ��P�����������P��zɯ��ξN�����!�F�x   x   r�s�(��uS����ƿ�Wݿ�O��������������O￧Wݿ��ƿtS��(��k�s�x�F��a �E��Jؾ���:���朾����朾1������JؾE��a �}�F�x   x   ��h� D��񀠿�R����ƿ��ӿ�ڿ�ڿ��ӿ��ƿ�R��􀠿D����h�T@�����E�D�۾O���ʢ���g���Ԟ��Ԟ��g��Ȣ��M���M�۾�E����T@�x   x   ��V��{���<��6��b����x��W���!6���<����{���V�P4�#S�S���Mؾz���T����������K����������T�t����Mؾ!S��&S�P4�x   x   ��?��z]���y�k�ʑ��z���z���ʑ�b��y��z]���?�w�#���
����ξ,��������������f碾l碾������������+��߄ξ�쾋�
�x�#�x   x   ��%�]j<�-Q���a���l�ӗp���l���a�-Q�]j<���%�;�����kK׾k���ί�����i�������碾1%���碾�����i������ί�k��lK׾���8��x   x   ˁ
�Y���)���3��H9��H9���3��)�K��ԁ
��6��7k־+��^���3��QU���霾�֞��L���碾�碾�L���֞��霾PU��'��`���(��?k־�6��x   x   ��߾/1��F��%|	����4|	�5��;1����߾{�Ⱦ�'��yk�����]��*���+���F����՞�������������՞�B���,���1���]�����vk���'����Ⱦx   x   %$�����`ž\�ʾN�ʾaž���$���"���<��P��P���E���C�)���m���	眾�f�����������f��眾o������D�@���U����O���<���"��x   x   }䂾�g��l
���b�g��o䂾�uw��j�t�b���a���h��uw�����ɱ���O���������h课	�������O��ӱ�������uw���h���a���b��j��uw�x   x   ��=���A��zD��zD���A��=��9���7��:���B��5R���h�{���$U�������į�-��������'���į�����"U��y���|�h��5R���B��:���7��9�x   x   �z�_g��+�Xg��z�Gl�l��E��,**��B�e�a������ ��N����[��+uξx>ؾ �۾x>ؾ,uξ�[��B���� ������c�a��B�-**�J�����>l�x   x   
5���}��b}��5��w���K+ڽv��������9��b�9B���Z��m	���5׾��쾎<��;�;��<������5׾}	��uZ��6B���b���9����5���c+ڽ����x   x   �+p��Ld�g,p��e��[s��~ ڽs��$�7�x�j��*������Q־����u�
��C����^S �����C�|�
������Q־����*��y�j�7�7����� ڽ s���e��x   x   �)+��)+�&�M�-]������[�Wv9�Tw������ȾQ�������#��<4�y@@���F���F�{@@��<4���#����V����Ⱦ���
Tw�2v9��[�(���K]����M�x   x   ���ò�d^V�ܩ��ǆ��,�*�n� מ���˾:���~K��"/��D��bT���^��Ob���^��bT��D��"/�}K�,�����˾מ�N�n���,�ņ�֩��^V����x   x   ���J�Т��(��L&/�_bx����xݾL��R,*��H�ic�z����3I��3I�����z�ic��H�[,*�X��xݾ���Abx�G&/�8������$�J�"��x   x   �TV�d������Q�0��g�N1��jj�����;��h`�Fn���d������oJ���ʥ�qJ�������d��Mn���h`���;����j�Z1���g�J�0����^����TV�
"7�x   x   [���I�콲�0�$���Щ���j���� �}oJ���u�K������<Z��jx���>ÿ�>ÿjx��@Z�����E����u��oJ��� ��j��˩��!�����0�V��d�����y���y�x   x   o��='/��i�Ū������]�%��S�͎��G6���Y��^dƿ��տܶ߿��޶߿��տ^dƿ�Y��I6��ˎ��u�S�d�%����������i�3'/�e��pǰ�I曽tǰ�x   x   ֽ,��ex� 4���m��g�%�SBW�l���g��������Lֿ������S ��S ��������Lֿ����g���k���YBW�b�%��m��4���ex�޽,�������ɽ��ɽ����x   x   b�n�����o쾎� �8�S�M���u4����ÿ^��Ĥ��F��J�����H��G��Ȥ��[����ÿy4��Q���0�S��� ��o����i�n�cI+�5r����0r�hI+�x   x   �۞�ݾ����tJ�U�������$�ÿ��M� �I����s��u�����F�M� ���&�ÿ|���S����tJ����ݾ�۞�$e�A�,�.��5��=�,�0e�x   x   �˾�����;���u�G:���ý�H��$� ��W�U��)"���$�("�V���W�"� �C�࿫ý�O:����u���;�����˾5f���7^���3�{�%���3��7^�6f��x   x   u���4*�Ur`��Ï�p_��YRֿ����"�Z��$�$���)���)�$�$�X��#�����XRֿj_���Ï�_r`�"4*�n���LX��ǋ�1]��<A��<A�1]�ǋ�RX��x   x   HS�$H��t��:����kƿN��Ɵ�w��K"��)���,��)�L"�v��ğ�Q���kƿ<����t��	$H�=S�{��h������h�c��V�c�c�����	h��m��x   x   -/�Wvc��l��.c��(�տ �����~��ѣ$��)��)�ϣ$������ ��$�տ0c���l��Vvc�-/��`��I̾��ZQ���Bs��Bs�YQ�����I̾�`�x   x   cD�z�r�����5�߿KY ��{��^"�V�$�a"�{���LY �;�߿���p�� z�aD����6,�a仾T]���Ɋ�*���Ɋ�S]��R仾@,����x   x   �qT����iU��$Kÿ��Z ����S��R��O��Q�����Z ���#KÿjU������qT��v'��C�v վ�a��mV����������nV���a��v վ�C��v'�x   x   ��^��S��ץ�YLÿ��߿�$��(����W]���%���$���߿ZLÿץ��S����^���2�r�n���^ƾ�w������������w���^ƾx��r���2�x   x   �bb��T��}W������}�տ�������� ��� �������z�տ����{W���T���bb�x�8�4������[־�>���ձ��ī��ī��ձ��>���[־ ��7��u�8�x   x   ��^��!��k���h��rsƿ�[ֿ����"俚���[ֿusƿ�h��k���!����^���8����)�e�ྰ�ʾ���ۄ��t���ڄ�������ʾd�ྺ)�����8�x   x   BwT�Qz�1r���Ȣ��h���ν���ÿ��ÿ�ν��h���Ȣ�3r��Kz�FwT�C�2�=���*�-E��Ѿbƾ�����P���P������]ƾ�Ѿ6E供*�9��C�2�x   x   @$D�ـc�m{��#̏�WD�����LA�����]D��%̏�i{��ۀc�=$D�S|'��u�$��X��3Ѿ"�Ⱦ�kž�Zľ-ľ�Zľ�kž%�Ⱦ-ѾV��$���u�Q|'�x   x   �6/�0H�M�`���u�����ٿ��޿��������u�N�`�0H��6/����H�A�꾊a־{�ʾ�ƾ�lž+�ƾ�Ǿ �Ǿ'�ƾ�lž�ƾ{�ʾ�a־;���H���x   x   �]��@*�� <�p�J�0	T�XW�3	T�j�J�� <��@*��]�i��8�S*վ{fƾ�D��������w\ľڈǾ�ȾۈǾ~\ľ�������D��~fƾT*վ�8�	i�x   x   (���>��(��)� ���%���%�-� �2��4��0���g��vW̾_﻾yj�����۱�M���T��!/ľ�Ǿ�Ǿ/ľT��Q����۱���|j��`﻾vW̾[��x   x   ��˾,�ݾL����� �����7��/�ݾ��˾�h���u��A���f��4^�����ɫ�v����S��K\ľ��ƾP\ľ�S��t����ɫ���4^���f��C���u���h��x   x   >ힾ/.���J��:õ�;õ��J��4.��DힾAu���Ӌ�HĆ�IZ��!ъ���� ���ȫ���������kž�kž��������ȫ�������"ъ�IZ��>Ć��Ӌ�Iu��x   x   ��n�؇x������Ď��x���n�^e�-N^��C]�@d�)Ps��/������	���ױ�*��kƾ��Ⱦvƾ(���ױ��	������/��-Ps�Ld��C]�N^�ae�x   x   ��,�8B/�0�0�M�0�3B/���,�+_+���,�X�3��IA���V�Ks�d̊��W���w��\=����ʾ"Ѿ Ѿ��ʾ`=���w���W��i̊� Ks�v�V��IA�]�3���,�_+�x   x   �����������^	��'�����W�%��CA��c�:R���\�� _��nZƾ~U־	��-;��྄U־pZƾ_���\��;R���c��CA�O�%����<��N	��x   x   ��������f������#᰽ ʽ<����Ţ3�=2]��������޻��վ��&��3"�6"�+���꾢վ�޻����x���:2]�ʢ3�����-ʽ'᰽x   x   xV���J�NxV���y�5���zʽ�v���,�6^�ċ��b���A̾!�W<�9i���|���;i�`<�� 쾫A̾�b��ċ�	6^���,��v��ʽ(�����y�x   x   �������67���y��ϰ�����NI+���d�b��kQ��/���Y�����k'���2��r8��r8���2��k'�����Y�2��hQ��'b����d�0I+������ϰ���y��67�x   x   �LݼB��<��؏��׽ϵ���W�x����^��2�����r�{i1��7@�G�I���L�C�I��7@�|i1��r���0���^��q�����W�ڵ�1�׽�؏�<�A��x   x   �����0��M���,ҽ4��JO]�����{5ž����&z��&2���J��^��/m�յt�ֵt��/m��^���J��&2�(z������5ž󢖾6O]�!���,ҽ�M����0�&��x   x   �<�>L����н;y���a�H����о���Ž%��E��zd����Ɖ�IE���}��JE���Ɖ����zd�#�E���%�����оO����a�;y���н<L���<�S8 �x   x   &ԏ�R+ҽay��c�9�{�ؾ�G���1���W�!�|�s��lҜ�����ֵ��Ե������oҜ�s���|���W���1��G�p�ؾ/��c�ky�W+ҽ9ԏ��^��^�x   x   ��׽t��e�a���#]۾G�ٝ9���d����Ri���������3Ŀ�!ǿ�3Ŀ������Ti�������d�͝9�G�1]۾��e�a�n����׽S���Q���P���x   x   ����Q]�K���őؾ�G��d<�U�k��i��?;��Ǿ��pͿHڿ��࿡��IڿpͿƾ��?;���i��W�k��d<��G���ؾP����Q]������㽓����������x   x   ��W�ť���о
J�!�9���k�����mm����Ŀ�fڿDG�����l�������EG뿏fڿ��Ŀim��������k��9�J��о������W�I��e;�� e�a;��L��x   x   [����:ž)����1���d��k���n���ǿL;Ῑ]�������������]��I;��ǿ�n���k����d�Ƴ1�'���:ža�����S���#�P��V����#���S�x   x   (d������Y�%�'�W���m>��e�Ŀ�<ῒ1��������8��������1���<�_�Ŀo>����%�W�P�%�����"d���`��8�S���/�<M$���/�1�S��`��x   x   k��I��	F�_�|�;n���û��jڿ�`�����'�l��m��'�����`���jڿ�û�7n��U�|�F�S��k������݅��B[��D��D��B[��݅�	���x   x   ��� /2�7�d��������vͿBM뿐�����[�����[��������?M뿛vͿ������>�d�/2����j;Ҿ����%���ۗk���`�ڗk�!���Ť��c;Ҿx   x   rz�|�J�_�ڜ�ʧ���ڿ����"����G��F����#�������ڿȧ��ڜ�X�|�J�}z�,�����ľ�ɡ�ތ��T���W���ތ���ɡ��ľ&���x   x   gs1�A�^��Ή�Ψ��j=Ŀ���ޥ�����f���)�i�����إ�����n=ĿϨ���Ή�B�^�es1����m㾙K��;椾����H������?椾�K���m���x   x   �C@�{?m��N��N���-ǿ�࿾�������������������	-ǿL����N��?m��C@�ow�����
׾�������������������	���	
׾����pw�x   x   �I�j�t�򇒿^����?Ŀ�ڿS�^h���:��dh��S뿎ڿ�?Ŀ^�������i�t��I�k�%�p2
����o�ҾK�¾����r'������L�¾p�Ҿ���r2
�h�%�x   x   :�L��t�rP��𫦿t����|Ϳ�rڿ�FῑF��rڿ�|Ϳt���񫦿oP����t�@�L�M+���������K!վ�L;EʾBʾ�L;I!վ�㾥�����M+�x   x   ñI�Dm�|҉�ߜ�"���˻�H�Ŀ_�ǿC�Ŀ�˻�$��ߜ�~҉�!Dm���I�>N+��x��q�S��Ɇ⾺kܾ��پxZپ��پ�kܾΆ�S���q��x�>N+�x   x   �H@���^�C����<v���G��qy��wy���G��6v����D���^��H@���%����r���򾕝�<G澶��]W�XW澱��9G澓�龇��r�����%�x   x   �z1��J�D�d�*�|�����u��Ǫ���u�����-�|�B�d��J��z1��|�,6
�����}����X��1U쾥�	��3U�[����}����-6
��|�x   x   ���92�IF��W��d��k��k��d��W�CF��92�
����K��������"��J澎V�p�Fy��By��l�V�J� �������J�����x   x   C�������%�k�1���9��w<���9�b�1���%����:��Q����y�׾��Ҿ(վ
qܾ���'�mz��z���nz��,ﾝ��qܾ(վ��Ҿ׾�y�U���x   x   3��-������X��W��W��X�	��!���4��*KҾ,�ľ�V��� ����¾�S;��پ�[�J�*{��.{��G��[澣�پ�S;��¾� ���V��&�ľKҾx   x   �u��MOža�о^�ؾvx۾a�ؾ\�оIOž�u��Xͬ�񱤾Pա�v�ũ��۲��zʾ�`پ\��r��\澌`پvʾڲ��ĩ��r�Uա�����Sͬ�x   x   X���ط��L���Q��^��J���ַ��e���o���酾���͖��Î��W����.���ʾ�پ����W��W�����پ�ʾ/��U���Ȏ��ʖ������酾
o��x   x   <�W��o]�b���c��
b��o]�*�W��S��S�'V[���k�����#P��������Q;roܾ{I�#�龀I�soܾ�Q;����죦�!P������թk�(V[���S� �S�x   x   ��� �������� ������J�#�a�/��+D�;�`�����0���A�����¾�#վ��⾶�龶�龀�⾆#վ��¾C���7�������%�`��+D�n�/�B�#����x   x   ��׽�Oҽ$�н�OҽV�׽ԧ㽡X��`���X$��&D���k�q����褾Q���1�Ҿ�㾖��������-�ҾP����褾n�����k��&D��X$�b���X��ʧ�x   x   a폽�e��te��w폽h���Ϻ��x⽦����/��G[������ɡ�J���׾X�������l��l� ���S�쾝׾J���ɡ�{���~G[���/����wx⽨Ϻ�J��x   x   A)<�x�0�5)<���^�㼍�?Ǻ�YF����#���S� ݅�n�����ľ�f�w���b,
�@�tp�=�a,
������f㾂�ľv���݅���S���#�uF��@Ǻ������^�x   x   ���'���K ���^���$��і���S��^��͹���4Ҿ_���O�6o���%��A+��A+���%�3o�K�i����4Ҿ˹���^����S�Ė��������^��K �x   x   ����c�ۼ7#��}��x��Ա��B��w��W��G@ξ���+��' �Y�-��
6��8��
6�W�-��' �,����M@ξ�V���w���B�ر�y���}�{#�f�ۼx   x   ��ۼH���2m��K��C=	�C��ф�>ҭ�Q:۾jr�v���w2�WTD��Q��W��W��Q�XTD��w2�r��fr�P:۾Lҭ��ф�xC�,=	��K���2m�����ۼx   x   �
#�h/m�kҵ�6~��D� J��f�����+��H�+��bF�v�]�sso��z�I�~��z�uso�r�]��bF�O�+�,��|��f��"J��*�D�:~�wҵ�o/m��
#�o�
�x   x   w�}��I��~�O�E� m���뺾kr����ؑ9�}~Y�{zv�/��������������/��}zv�v~Y�ґ9���vr��뺾m��F�E�~��I����}���E�БE�x   x   t���<	���D��m��^＾���g'�5D�(Si�y3��oc�����v}�����x}�����nc��z3��0Si�2D�_'����e＾�m����D��<	� t������v�������x   x   7��;C�^K�������UY!���I���s�	X��<ՠ�����Ⱥ��]���]���Ⱥ����:ՠ�X����s���I�XY!�׀����\K��8C�C��oнM歽G歽oнx   x   �B�|ӄ��h��v�2)���I�kw�����mB��$麿7Iɿ�Wҿfoտ�Wҿ7Iɿ&麿pB������kw���I�4)�v��h��{ӄ��B����H�ٽH뽧��x   x   �x���խ����B���D���s�|����ժ�!��� �ҿ�X߿I��K�忍X߿��ҿ����ժ������s��D�@����辎խ��x���|D����
��
����|D�x   x   �Y���?۾X���9��Xi��Z���D��X�����տ�+�6~�!��3~��+濎�տW����D���Z���Xi��9�Y���?۾�Y��(��)M�k90��&�m90�)M�(��x   x   (Eξ�v�`�+��Y��7��;٠��캿��ҿ?-���G]��H]����;-濧�ҿ�캿<٠��7���Y�`�+��v�,Eξ[��Vk�� �^��qL��qL��^�Vk��[��x   x   M������jF�k�v��h��%	��@Nɿ�\߿3���^��F���^��6��\߿>Nɿ$	���h��q�v��jF����J��X�ľn����ቾ|)z���q��)z��ቾw���Z�ľx   x   y��2��]�R5���!���Ϻ��^ҿ��忥	��[`��Z`���	�� �忈^ҿ�Ϻ��!��Q5���]��2��-���|��5�������Ϗ�Ϗ�����0����|��.��x   x   �. �y^D�c�o���������e��Swտd����~"��!��d��Owտ�e���������i�o�y^D��. �t����޾ZKþS��:U��䊦�8U��S��\Kþ��޾w��x   x   �-��'Q�0�z����4��g��aҿ�`߿�2��2��`߿aҿg��5�����)�z��'Q��-��l�����޾�;��þP���T�����þ�;�޾����l�x   x   �6���W�5�~��������Ӻ�/Sɿ�ҿt�տ�ҿ-SɿӺ��������>�~���W��6�~"�k�y������Z�ܾ��ؾ��׾��ؾc�ܾ���w���k�~"�x   x   �9�F�W�d�z�ӷ���%������󺿵��������󺿛���%��Է��^�z�C�W��9�F7 �5(�s�����N��O��S��P��G��M�����s�2(�F7 �x   x   =6��+Q���o��9���n��Q࠿M��bߪ� M��T࠿�n���9����o��+Q�>6�Y8 ��y�=��n���� �2�A%�R��F%�	2��� �o��>���y�W8 �x   x   ��-��dD���]���v�l>���b��ڸ��߸���b��i>����v���]��dD���-��%�*�%��`���1-���	�!p�p���	�3-���`�$��*��%�x   x   f5 �T�2�juF���Y��gi�4�s�E~w�1�s��gi���Y�nuF�S�2�c5 ��q��n��u�'������?	�����D�|���D�����?	����(���u��n��q�x   x   4����+���9�>%D�%�I��I�?%D���9���+��8�����������+���� ��.�����M�aR�^R��M�����.�� �/�������������x   x   "'���������#8�~i!�-8��������'��]�羬�޾޾�����B5�[�	�nF�2S���2S�pF�Z�	�E5�����޾��޾_��x   x   (Vξ�S۾��
������������辈S۾&Vξ!�ľމ��WþQ;!�ܾ��)�Cs�Ѓ��S��S�σ�As�)���,�ܾP;Wþ׉���ľx   x   �i���签}�������z��}���签�i���i��~��P���w^��{�þ�ؾšﾂ���s�wG��O�sG��s��������ؾy�þz^��T������zi��x   x   ���sㄾ�\���������\��lㄾ+���b���w��J퉾���1`�������׾���p)�M�	�x��z��P�	�j)����+�׾����3`�����C퉾�w��d��x   x   d0B��4C�E�o�E�	E��4C�c0B�œD��>M��^�>z�@ُ����2���=�ؾ��ﾫ5�0��A	�0��5����3�ؾ.������@ُ�>z��^��>M�ГD�x   x   ��� R	�����R	�������(�K0�Y�L�r��׏��]��ϵþ٤ܾ����� ��������� ����ڤܾҵþ�]���׏��r�S�L� K0��(���x   x   ���.j��u�1j������z�н;e뽚(
���&��L�*7z�1��EY��;���z��������{������	;@Y��,��;7z��L���&��(
�<e�v�нx   x   n�}�>\m�W\m���}�w���W���G ٽ�$
�AC0�c�^��剾ڃ��Nþ޾4���r�=��<��r�<���޾	Nþユ��剾Z�^�HC0��$
�Z ٽJ���M���x   x   �(#�m���(#�ѰE����4����U���f.M�Vm�������|����޾���h� $��t�$� h������޾�|������Ym��c.M����U�,���5��ӰE�x   x   ��ۼ�ۼ��
�^�E�T����wн$���~D�B���Y��b�ľ�群���g���r/ �p/ ����g������]�ľ�Y��E���~D�*���wн3���5�E�n�
�x   x   �d��J���)��`�W����}���x/���j������L��c�P���l�t���B%��'��B%�s���l�N��cྲL������}�j��x/��}��u����`�(*�J��x   x   �>��޺��DM�⽠��g�7+��Di�y����t��@�#�	�̟�1P,���7�]f=�af=���7�/P,�П�&�	�@꾽t�������Di��7+��g�۽��mDM�����>��x   x   ) ��@M�~A��R�뽥�)��j�������Ǿ�����k��2*�v>�Y�M�[TW�a�Z�XTW�_�M�t>��2*��k�������Ǿ�����j���)�W�뽛A���@M�G �9�x   x   �`�뺠�q�뽧�)��\l�����awξ\���	�"8�R�P�� e�[{s�� {�� {�Z{s�� e�W�P�"8��	�[��kwξ�����\l���)�[��ຠ��`�5O0�jO0�x   x   �����d�i�)�=]l�_ ���pҾ�����$�6�C���a��6{������ƍ��鏿�ƍ������6{���a�;�C���$�����pҾ_ ��D]l�p�)��d����f��_�m�X��x   x   7w���6+���j������qҾ�p�\�(��	L��Yn��������<���2L��1L��<�����~����Yn��	L�a�(��p��qҾ������j��6+�Aw��n:��⤽	⤽y:��x   x   !v/�Ei�H����yξ���F�(�z�N��?u�񶌿�`���r�����%�������r���`�������?u�u�N�C�(�����yξF���Ei�v/�\�r���սq��\�x   x   ѫj�������Ǿ���?�$��L�Au�͎�W��g��Ὼ��C���C��⿺�g��T��͎�Au��L�?�$������Ǿ����ҫj��E9��B�^�^��B��E9�x   x   �����w�����t�{D��]n�����V�������_��7�ȿV�˿5�ȿ�_������V�������]n�zD�w�����w������_�r�sK�m5��U.�"m5��sK�^�r�x   x   �M���D꾦o��8��a�����ic�����a����˿��ѿ��ѿ��˿ a�����jc�������a��8��o��D��M��\0��
���0h��[��[��0h���R0��x   x   f���	��8*�ݳP�J?{�,����v��Tú���ȿ�ѿ6	տ�ѿ��ȿTú��v��*���J?{��P��8*���	�'f�Aպ����,��l���,�� ��Iպ�x   x   �����.>�U
e����᝜����H���˿d�ѿc�ѿ�˿�H��!��᝜�!���P
e�)>�������(ܾ��������楾v���s����楾��������(ܾx   x   �p�W,���M�$�s��͍��R�������I���ȿJ�˿�ȿ�I�������R���͍�'�s� �M�W,��p������k߾�cξ��ľD��|ﾾD����ľ�cξ�k߾����x   x   ����7��_W��{�C��S��E���ƺ��e���e���ƺ�F���S��E񏿏{��_W�	�7�����,
��E��W����Wp߾�`޾�`޾Rp߾���_�꾬E��,
�x   x   %I%�Vp=�Z�Z�&{�Iύ�Ǡ���z��� ��RŲ�� ���z��Ƞ��Fύ�${�a�Z�Xp=�)I%��Z�����?��Z��5����k������k��C����Z���?�����Z�x   x   ��'��q=��bW�Ƌs�����ȍ��@i��V��Z��Ai��ō������ʋs��bW��q=���'��'�Y���	�� 	���
�w����r����
�� 	���	�Y��'�x   x   VK%���7�P�M��e��H{��Æ�ȿ��7Վ�ÿ���Æ��H{��e�S�M���7�YK%��(����H�����������
�<��
�����������H����(�x   x   ���\,��&>�Z�P���a��kn��Pu��Pu��kn���a�Z�P��&>��\,����]��Z��I�q�XH�v����$�C�'�<�'���$�{��WH�n��I��Z��]�x   x   \v�`���A*�� 8�ND�xL��N�{L�HD�� 8��A*�_��Zv�'1
�F��R�	����XI�{!���)�+9/�X51�39/���)�{!�ZI����O�	�E��'1
�x   x   ���:�	��y���O�$��	)��	)�O�$���|y�8�	����m����O���C��$	�j����ˣ)���1�=H6�9H6���1�ͣ)���j���$	��C��O��j���x   x   hu�jV������`��6~�g�������nV�mu�F6ܾx߾Z���d���
����ӗ$�R;/�RI6���8�RI6�T;/�ӗ$�����
��d��]��x߾F6ܾx   x   r]��������Ǿ��ξ0�Ҿ-�Ҿ��ξ��Ǿ����m]��\㺾=���Cpξ��⾙���ʵ���M�'�r81�BJ6�FJ6�q81�I�'���˵��������=pξ9���a㺾x   x   �������s��
���3���	������������#>��Q)��~�����ľ}߾!x���|A���'��</�T�1��</���'��A��x��}߾��ľ����P)��>��x   x   =�j� ai�r�j�|l�&|l�h�j�ai�J�j�Ĩr��+������k�#Q���m޾-���_�����$���)�æ)���$���]�;����m޾!Q��e󥾒����+����r�x   x   Ќ/�:N+���)�A�)���)�6N+�ٌ/��[9���K��Gh��8��ߗ��V����m޾x�����x��5��~!�/�x�����vx���m޾Y���ޗ���8���Gh���K��[9�x   x   �������`�D콦�𽇜���n�WU���5�$[��v�������O��M|߾ۦ���
�3��)L�-L�7���
�ئ��P|߾�O�� ����v��[���5�NU��n�x   x   ���~נ�;]��yנ�����W��X�㽨m�?f.�q[�g6������ľ���d���$	����� �����$	��c�������ľ��e6��p[�Jf.��m�Q�㽮W��x   x   �;`�ShM��hM��;`�0'�������%ս�j��z5�T?h���������jξ���8B�\�	��I��I�\�	�?B�����jξ�������Q?h��z5��j��%ս����'��x   x   �;����|;�m0�n������K�7}K��#��� ��)���o߾\G�����X����X����VG��o߾.���� ���#��9}K��K��㽳�gn�m0�x   x   rY���Y���*�\c0�0���E���a�RK9���r�]2��eֺ��(ܾ����u*
�fW��#��#�hW�z*
������(ܾcֺ�`2����r�]K9��a��E��%��-c0�O*�x   x   ƀ��#�����cVH�����O��� �>�W�~��=���D�ξ�i�J�����!���!���H���i�F�ξD�����7�W��� �O彑���SVH������#��x   x   ���ˮ߼U�2������<ӽ���ѡM�Ú�����P�ξ_��@
�K��^�!���&���&�[�!�I��C
�i��F�ξ���˚��סM�����<ӽ����-�2�y�߼|��x   x   w���2�-��TH˽���ZI�l��������Ҿ����3�g,"��_/��7�q�:��7��_/�g,"��3����.�Ҿ����c����ZI���TH˽C����2�gw���VӼx   x   �HH������F˽k���H��Ѕ��&��e�ؾ�9�����N.�JW?��K���Q���Q��K�FW?��N.�����9�]�ؾ�&���Ѕ��H�q���F˽����qHH�� �� �x   x   ��7ӽ��LH���������ݾ�@�!��:�?QO��_��1j���m��1j��_�>QO��:�C�!���ݾ�������NH����7ӽ����#Mv�la�Mv�x   x   �D�����YI��Ѕ�����{߾��
��J'��VC���\�;�q������e���e������>�q���\��VC��J'���
��z߾�����Ѕ��YI�����D���j���r�����x   x   -� ��M�_����'��c�ݾ�
�N)�oH���e�ѱ��ɉ�����2������ɉ�ϱ���e�oH�N)��
�j�ݾ�'��^����M�*� ����Z�⽵r׽R�⽚��x   x   M�W�����k���νؾ���L'�.pH�.i�w���P؏�)���?&��>&��*���R؏�v���.i�.pH��L'���ýؾi�������I�W���2����{��{�������2�x   x   �	��̺��k�Ҿ<�,�!��YC�9�e�?����L���,�������,��K���@���<�e��YC�(�!�<�v�Ҿͺ���	���k�_OO���?�.;���?�bOO��k�x   x   ڤ��L�ξ4���J��z:���\�J��ڏ�@ ��꘦���똦�@ ��
ڏ�I����\�|:�J��1���?�ξۤ��]є��F��gNx�^�o�X�o�^Nx��F��Vє�x   x   ��ξ��7��S.��WO�r��̉�흘��.������H	�������.��흘��̉�r��WO��S.�7�����ξJ���pg���ٛ������������ٛ�sg��R���x   x   �iﾭ

�41"�^?�C�_� ���-��*����������������*��,�����G�_�^?�21"��

��i��־-ƾ
Z�����y��y�����Z�� -ƾ�־x   x   !������e/�<�K��;j�k��8���*���0��󛦿�0�� +��8��k���;j�=�K��e/����!�����d�B�޾�)ܾ��۾��۾��۾�)ܾJ�޾�d徼��x   x   {�H�!���7���Q�j�m��k���������$��$����������k��p�m���Q���7�D�!�x�o(�.` �b�������, �����, �����h���1` �k(�x   x   �$���&���:�F�Q��>j�f���gЉ�~ޏ�{���|ޏ�iЉ�h����>j�E�Q���:���&��$������n+���W����������]���j+������x   x   đ���&��7�!�K���_��r��������������r���_�#�K��7���&�������,���J�^e�6Z�s$�	\'�
\'�s$�5Z�be��J�)�����x   x   �&�q�!��j/�;d?�~_O���\��	f�3;i��	f���\�~_O�;d?��j/�p�!��&�����-����� �?�)�~�1�-<7��79�2<7��1�;�)��� ����-����x   x   R�����7"��[.� :�
eC��|H��|H�
eC� :��[.��7"����O�� �����Xe#�e/�"3:�S�B�`�G�X�G�O�B�'3:�e/�Ue#������ �x   x   {��
��>�`����!�fX'��Z)�kX'���!�^���>�
�|���,����M��� ��/��$=���H���P�ӲS���P���H��$=��/��� ��M����,�x   x   sv���������E�y���
���
�z��E��������mv�3��Se �0�hi���)��5:�I�a(T��'Z��'Z�_(T�I��5:���)�ii�0�Qe �2��x   x   ��ξ��ξ}�Ҿ��ؾòݾ��߾ǲݾ��ؾx�Ҿ��ξ��ξ
־�p�. �����i_��1��B�[�P��(Z�a]��(Z�\�P��B��1�g_����0 ��q�־x   x   %����ɩ��Ǫ�@9��H
��K
��>9���Ǫ��ɩ��������:ƾ��޾`���� �py$�B7�i�G�ǶS�C*Z�G*Z�ȶS�e�G�B7�ry$�� �]�����޾�:ƾ���x   x   =��˧������&���O%��#������ħ��:���ޔ�u��h��X8ܾ�3 �Y��Wc'��>9�f�G���P�	,T���P�i�G��>9�Uc'�V��3 �^8ܾh��u���ޔ�x   x   ��W�ϷM��rI��!H��!H��rI�ϷM���W��*k��S���盾}%��7�۾�%�����c'��C7���B�JI�PI���B��C7��c'�����%�6�۾x%���盾�S���*k�x   x   A� ����d����n����H� �j�2��fO��gx����懷�Lܾ�%�)��,{$�
�1��9:�d*=��9:�	�1�2{$�'���%�Lܾ凷�����gx��fO�n�2�x   x   �g�&Yӽ(g˽g˽-Yӽ�g�̯����@��p�W�������C�۾4 �O"��a�6�)�r/�u/�;�)��a�L"�4 �C�۾����\���}p��@�}��ͯ�x   x   î��Ό��"���͌�̮���7������� ;��p�W��`$���7ܾ?������k�v� �j#�t� ��k���H����7ܾ]$��Q���p�" ;�	����⽿7��x   x   SoH��2��2�LoH��wv�Š�~�׽���n@�0bx��䛾�e���޾�����0��O������O��0�������޾�e���䛾2bx�k@������׽Š��wv�x   x   ݩ����߼����� ��'a�����X�⽐���]O��N���o���5ƾ�l��c ���Y��/�^�����c ��l得5ƾ�o���N���]O����a��w����'a��� �x   x   !1��1��0xӼٔ ��ev��)�����2�ck��֔������־]��)���ޚ�ٚ����)�^��־�����֔�\k�"�2����)��fv��� ��wӼx   x   ��a��0��%�߼�7�_��W�ս�����J��:���G�¾�x��"��!o�J�C�N�!o��"���x�I�¾=������J����^�սJ��Ӷ7�3�߼�0��x   x   �%��|TƼ�� z�o���k��7��p�a���2���o�ؾ������sL�f��d��qL�������s�ؾ-���^����p���7��k����
z���zTƼ�%��x   x   ȵ߼�z��n��Q�����Y@-��He�^��>����R׾ij��r�
����{�h��|����q�
�cj���R׾F���^���He�\@-����Q���n��z���߼���x   x   ͦ7��
z�'O��������(�@g`�W}���K����پ ��������)�(�D.�E.�)�(�����������پ�K��V}��@g`���(�����#O���
z���7��"��"�x   x   g������y����(��_�] ���a����ݾ���yL�ۏ(���5��>��jA��>���5�ڏ(�vL������ݾ�a��] ���_���(�v������p��}�l�65\�h�l�x   x   +�ս�f�s=-�f`�T ��	����{����:��1��B��N��
U��
U��N��B��1�:�����{����W ��f`�r=-��f�#�ս����0���A��� ���x   x   ғ��7��Ee��|��b��&|ྺ���l �p�7�\bL��Z\��wf�:�i��wf��Z\�ZbL�p�7��l ����$|�b���|���Ee��7�ӓ�� ���轃�ཱི��� �x   x   ��J���p��\��L��j�ݾ���Mm ��:��Q�?je��zs�^�z�\�z��zs�Bje��Q��:�Lm ����m�ݾL���\����p���J��01�9�!��o��o�@�!��01�x   x   ꂾ�������2�پN��5�E�7�<�Q�_�h��lz�
߂�τ�߂��lz�]�h�>�Q�G�7�4�L��2�پ�������ꂾ�i��X�`�O���L�d�O��X� �i�x   x   *���T���S׾H��3O�f�1��eL��le�Nnz�ZĄ�x���w���[Ą�Rnz��le��eL�g�1�4O�J��S׾K���(����V��Iǋ��;��zU��xU���;��Lǋ��V��x   x   [�¾r�ؾ`l��c���(�ИB��_\�s�����K���n���K�������s��_\�ΘB��(�c��\l��w�ؾf�¾P����B������ب�����B��좭�V��x   x   ;s����j�
����q6�j�N�~f�B�z�pф�������qф�A�z�~f�k�N�u6����k�
����2sᾴCվ�Ͼ��ξ�ϾO�оM�о�Ͼ��ξ
�Ͼ�Cվx   x   ���������x�(�އ>��U�:�i���z�4₿�Ƅ�2₿��z�?�i��U�ڇ>�w�(����������:���n�t�u��=������=���u��x��n�9��x   x   �m��M����.�sA��U���f���s�rtz�xtz���s��f��U�sA��.����M��m��h��d���	�r��i��S
�T
�i��o����	��d��h�x   x   ���������.�E�>�N�N�e\��se��h��se�	e\�O�N�C�>��.���������`�Um����0�I$&��+���,��+�L$&��0���Vm�a�x   x   rC��������(�6���B�JmL�`�Q�a�Q�JmL���B�6���(������mC�����p�N�!��1,�6�P�>��
C��
C�M�>�6��1,�M�!��p����x   x   ���P�������d�(�P�1���7�R":���7�O�1�c�(��������P���~��#��8�&�W4� UB�(N��V���X��V�)N��TB�W4�:�&�!��~��x   x   Vq���ض
�����V�;$�fw �bw �:$� W����ٶ
���Rq�*��r�N�&�[7���H�?X���c��Bj��Bj���c�CX���H�[7�P�&��r�)�x   x   �(��P���py��K$��ў�]��� �`��Ξ�I$��qy��K����(��@m�%q�y�!���4��H�5�[�U<k�u�u�K3y�z�u�R<k�4�[��H���4�x�!�&q�>m�x   x   Iᾄ پ_a׾��پ��ݾ��ྈ�ྟ�ݾ��پba׾� پDᾇ��j���"6,��XB�X��=k�W�y���������V�y��=k�X��XB�"6,���j����x   x   ��¾���	���[��dr�����ar���[����������¾�Pվ�{��
�/7���6��"N�M�c���u�����4���������u�N�c��"N���6�07��
��{�Pվx   x   ���������j��=����.���.��<����j�����������+��"�Ͼ����+&���>��V�Ij�)8y�\���]���+8y�Ij��V���>��+&����#�Ͼ,��x   x   ������p��^e�.`�r6_�1`��^e���p����zd��J���Ͼ������s+��C�B�X�iJj���u��y���u�jJj�D�X��C�r+�������ϾF���vd��x   x   ��J�<�7�S-���(���(� S-�E�7���J�5j�Ջ�R����Ͼ�N����H�,��C�*V�-�c�oCk�tCk�0�c�'V��C�H�,����N����ϾR��
Ջ�8j�x   x   ݧ��y��0��*���0���y�ܧ��F1���X��I���&����оb���G��+�p�>��&N��"X���[��"X��&N�s�>��+�F�^�����о�&���I����X��F1�x   x   ��ս����j���j�������ս:� �=�!���O�~c���訾��оP��b��o.&���6�N^B��H��H�Q^B��6�l.&�b��P����о�訾}c����O�A�!�2� �x   x   ���8z��.n��7z�����Ȳ�o��r��+�L�c��U&���ϾЇ��ע�S:��:,���4�Rb7���4��:,�T:�ڢ�̇��	�ϾU&��c��)�L�o��w���Ȳ�x   x   D�7�%��2��1�7�=m��ס������U�O��H��FQ��:Ͼ���
�����!�γ&�γ&���!����
���=ϾGQ���H��Y�O�����རס�bm�x   x   ��߼yƼ��߼�?��X\�.ԡ���轤�!�x�X�oҋ�1����Ͼ&|�7k�Hs��u�m���u�Hs�4k�(|��Ͼ/���qҋ�s�X���!����'ԡ��X\��?�x   x   �<��~<��M)��9�,m�6���1� �J>1��i��_���'��:MվO���l����������l�T��7Mվ�'���_���i�Q>1�)� �1���em�9�1)��x   x   RmT��C��-�Ӽհ.�������̽���@�C�:}�CG��qX��K�پh1�|�U�	����W�	�|�a1�I�پvX��DG��4}�=�C�����̽����԰.���Ӽ�C��x   x   �8��eS���v�<d��'��5���^M'�Gq[��z��R��F�ž�྘���[l�����Yl�������D�žN���z��Kq[�YM'�'���(��Ld��v��S��z8��x   x   �Ӽ�p��U��~���xܽ2���0G��}�3}���}��P׾��ﾞ��H��G�	�K��������Q׾�}��4}����}� 1G�7���xܽ�~��qU��p���Ӽ⹼x   x   7�.��
d�Z{��s�Խ�}���<��q��L���>����Ӿc��g��1���Y��Y�1��h��d����Ӿ�>��L���q���<��}�q�Խa{���
d�)�.���ȉ�x   x   ������Prܽx|���9���l�繓�������Ծw�������<{����<{�������s�󾏈Ծ����鹓���l���9�v|�Orܽ�������=l�q�_��=l�x   x   ��̽���c����<���l�:�������R־����������#�{�(�~�(���#���� ������R־����7����l���<�f�������̽0⳽GZ)⳽x   x   ���=D'��*G���q�P���Ŗ��A,׾5S��c%�
 �V�,�s4��+7� s4�Y�,�	 �_%�8S��B,׾Ɩ��P�����q��*G�=D'�����d�����������d�x   x   ��C�Df[���}��J��F����S־�S���|�Ո#���2��=�HZC�GZC��=���2�؈#��|��S���S־H����J����}�Cf[���C�(R4�d�+�=�'�;�'�l�+�(R4�x   x   ��|��t���y��r=��=�Ծn	��x&���#��4��B��fK��jN��fK��B�	�4���#�w&�p	��=�Ծo=���y���t����|���n���f��sc��b��sc���f���n�x   x   �=���x��.z��o�Ӿ������ ���2��B��6N�MT�	MT��6N��B���2� ������r�Ӿ1z���x���=��Ea��������蔾蔾
������Aa��x   x   KN����ž� ׾k�ﾭ�������,��=�iK�JNT�aW�JNT�iK��=���,�������k�ﾾ ׾��žPN��h���Z$���_������m������_��X$��j���x   x   �پE�྘��ǡ�����#��w4��^C�/nN��OT��OT�3nN��^C�w4��#����ɡ����D���پeCپtlݾ>���=�r��u���=�=��xlݾdCپx   x   �'�����������Y���(�M17��_C��kK��:N�kK��_C�P17���(�Z������������'�~������ml���
�_�����_����
�ll���������x   x   �w��j�C��0]����͐(��y4���=�֦B�ܦB���=��y4�̐(����1]�G���j��w�����AQ�\���&�3*�3*��&�]��CQ�����x   x   ��	�6��'�	�^�J��"�#��,��2���4��2��,�"�#�L��^�$�	�5����	�ME�>��,&�KB2�X�<�ӖC�|F�ԖC�W�<�JB2��,&�>�ME�x   x   �������8�n����� ���#���#� ����n��7��������,����!���0��@�J3O�5Z��'`��'`�5Z�K3O��@���0���!�-��x   x   t�	�:m��������(���-�ۄ��-�&���������;m�v�	�!���$��j6��I���\�z#l��`v���y��`v�y#l���\��I��j6��$�!��x   x   {�� �����E�������^c��Zc�������D������ ��{�H���!�l6��-M�S�c��w��O���P���P���O���w�R�c��-M�l6���!�H�x   x   A1���
׾��ӾǖԾ6b־�;׾8b־ȖԾ��Ӿ׾���J1�~��B��0�� J�ӿc���{�1������L@�����1�����{�Կc�� J��0�B�|��x   x   ��پ��ž����fJ��鿳�䤳�椳�迳�cJ��������ž��پ����{��2&�#�@��\�b�w�����W�����������W�����a�w��\�#�@�2&�|������x   x   [��J������zW��,Ɠ�!��+Ɠ�}W�����H���[��{Pپd���,X�CI2�:O��)l��R������ ���m��� �����R���)l�:O�DI2�,X�]���{Pپx   x   �J�� ��	~�$�q���l���l�!�q��	~�《��J��Kȸ�Q{ݾXt�����<��=Z��hv�kT��5C��������5C��kT���hv��=Z��<����[t�Q{ݾJȸ�x   x   �}�J}[�l@G�k�<�7�9�s�<�g@G�D}[��}�o���3�������
�D�&���C�2`���y�FU��V���Z��V��FU����y�2`���C�D�&���
��㾗3��o��x   x   2�C��X'��������������X'�5�C�B�n�E,��jp��\P龉���=*��F�a3`��kv�U����������U���kv�b3`��F��=*����\P�cp��K,��M�n�x   x   #��!�����ܽ��ԽĐܽ+������h4�)g��˔�՟��_��}���>*� �C�?AZ�7/l�Һw��{�кw�9/l�?AZ� �C��>*�{��a��۟���˔�g��h4�x   x   Z�̽)9��������9��P�̽�w��+�8�c����4����쾦����&���<��?O�*�\���c���c�*�\��?O���<���&������,������B�c�#�+��w�x   x   r���~3d��:U��3d���������������'�a�b�.�������[R���
����N2���@��J��7M��J���@�N2������
�[R龏���0���T�b���'���������x   x   >�.����Ќ�1�.��il��	��`����'�g�c��˔�uq����㾻v��[�.7&���0�t6�t6���0�-7&��[��v����oq���˔�o�c���'�N���	���il�x   x   mԼzt���Լ���*�_����V�����+���f��+��L4���}ݾ˱�����F���!�� $���!��F���ȱ���}ݾO4���+����f���+�a�������_����x   x   mN��JN������_l�J���@s�d4��n�}m���Ǹ�yQپ�������K��������K�������zQپ�Ǹ�|m���n�d4�8s�L���$_l�!��>��x   x   ��Y�Y-����Ӽ��,�:̇��Nʽ;�:�A���z�粛��N�� ׾�>����h�	���>���׾�N��粛���z�8�A�;��Nʽ,̇���,�
�ӼO-��x   x   �!��x��^��7W�g��A���o�bQM�㝁����8+��Ҿ9��>d��~��{��:d��=�� Ҿ3+�����杁�gQM��o�.��g���7W�'^��x���!��x   x   d�Ӽ)W��+E�ܺ���Ž�	��v0�,�`��W�������Խ�.�Ӿ���ﾊ<�����(�Ӿ�Խ������W��'�`��v0��	��Ž⺌�i+E�W��Ӽ ���x   x   ��,��(W�۶�����^��~� ��L��C}�'Q��c���,ɾ��ܾ|�3��0��|꾵�ܾ,ɾd���&Q���C}��L�|� ��^��l��嶌��(W���,��M��M�x   x   ���{Z��ŽsZ��R�"�C�nMq��Ñ�򰫾T�ľۧھ��뾽��������������ܧھT�ľﰫ��Ñ�lMq�&�C�L�uZ��&ŽoZ������is��Uj�js�x   x   �7ʽ����^� �S�C��m�H��aK����þ�JܾN����������������K���Jܾ��þbK��K���m�V�C�a� ������7ʽQ���~���~��A��x   x   ,��c��m0�)�L�WJq����������þʨ޾���Y���
�l���
�[�����Ǩ޾��þ�������XJq�(�L��m0��c�,�}<��%�����%��<�x   x   FA� BM��`��<}������J���þk�߾G��-J�7x�������7x�,J�I��k�߾�þ�J�������<}���`�$BM�KA��M;���8�]�7�[�7���8��M;�x   x   Srz�𔁾�Q��UM��S�����þ��޾���	�����0�9p��0�����	�����޾��þR���QM���Q��򔁾Lrz�U�w���x��6z��z��6z���x�[�w�x   x   ���%���Ѻ������_�ľ�Kܾ���>K������� �� ������<K�!����Kܾ\�ľƻ��Ӻ��#�������?,���p��.�����������3����p��;,��x   x   �@��� ��Pν�-ɾ��ھ���,��#z�X2�b� �O�"�a� �U2�%z�-�������ھ,ɾLν�� ���@��E�����ƾ�ξ9Ӿ�վ9Ӿ�ξ��ƾE���x   x   �	׾�Ҿ�Ӿ��ܾw��������
�����r�S� �T� ��r������
�����v����ܾ�Ӿ�Ҿ�	׾��ྩc�A������Ɯ�Ȝ����?����c���x   x   ���R��ٹ�g{�������������24���/4�������������c{�ֹ�U�澀�ﾷ��'���9�RY������!����SY��9�&�����x   x   ;��R[������P��������
��|�.��0���|���
����I�������O[��9������}���%�(�1�M�:�՟?�ӟ?�M�:�,�1���%��}����x   x   �������::�����������t��YO���	�WO�r�������������5:������������$�Z�5���E��yS�5i\�ŉ_�9i\��yS���E�\�5���$���x   x   ��	�� ��(����m��6��(���h"��h"��+���8��m����)�ﾉ ����	�~o�{k,��BA���U�"Rh�*v��o}��o}�,v�&Rh���U��BA�{k,�o�x   x   M��`�����͏ܾG�ھ�UܾE�޾۾߾D�޾�UܾH�ھ͏ܾ���`��M��wp��/��OG��8`��pw��6���r��m����r���6���pw��8`��OG��/�wp�x   x   ���Ǵ�K�Ӿ5ɾG�ľj�þf�þg�þl�þE�ľ4ɾR�ӾǴ澌������m,��PG�#�c�Jf�ǋ���	��������ǋ�Hf�#�c��PG��m,����x   x   ��NҾ8ؽ�Ʊ�	����U���Ĩ��U��
���Ʊ�4ؽ�HҾ����˲$�{FA�s;`��g�^������nL��9�jL������`���g�r;`�{FA�̲$���x   x   �׾�+���Ť�X���̑�`#��`#���̑�X���Ť��+���׾S$��̓�3�5�} V�iuw��ȋ����������v���v�����������ȋ�iuw�~ V�2�5�̓�Y$��x   x   M��մ���\���Q}�w^q���m�z^q��Q}��\��״��M�����I��+�%�6F��Yh�e:���Ŕ��N���w��|M���w���N���Ŕ�e:���Yh�6F�+�%�G�� ��x   x   ܲ�������`���L�*�C�)�C���L�	�`�����ڲ������is�oB�^�1�1�S��v��w��6�������y��y������8����w���v�0�S�_�1�qB�gs����x   x   �z��WM���0�C� �F�G� ���0��WM��z�|:����ƾv���ac�4�:��t\��{}����?����P��K����P��>�������{}��t\�5�:�^c�y�����ƾv:��x   x   ǕA��v�T��v���v��R��v�ΕA��w�W����!ξ�����3�?�Ӗ_�@}}�Uy���Ȕ����������Ȕ�Vy��C}}�Ӗ_�2�?�������!ξ[����w�x   x   b?���佪,Ž����,Ž���`?�ce;�;�x�5ϣ��LӾ���=�!�@�?�Nw\�lv��=��_͋����_͋��=��jv�Kw\�A�?�<�!�����LӾ5ϣ�/�x�be;�x   x   VWʽ�s��Uˌ�Yˌ��s��YWʽ2P�?�8��Tz��ӥ��,վ������5�:���S��`h�e~w��r��r�d~w��`h���S�7�:��������,վ�ӥ��Tz�C�8�6P�x   x   ԇ�VNW��HE�vNW�ԇ�K-���9���7�{�3ԥ�aNӾ���Nf��1��F��V��E`��c��E`��V��F��1�Jf����kNӾ5ԥ�{���7��9�C-��x   x   ��,�	q��p���,���s�����a��b�7�EUz�jУ�i$ξI���2F���%�L�5�MOA�5[G�7[G�NOA�J�5���%�6F�N���a$ξfУ�JUz�i�7�^��Ҝ����s�x   x   o�Ӽa���ĮӼ�l��j�B����8���8�׽x�ց����ƾ�x�K��E��̹$�v,�5/�v,�ʹ$�G��K���x���ƾف��׽x���8��8�J����j��l�x   x   7��7��?���>h���s�h(���M��c;���w��;��[�����ྒ+�������w��w������+�����Z����;����w��c;��M�q(����s�dh�����x   x   ��o�D����Mݼ�R1����|�̽���wC���|�����Y���YPؾ�!�}#�.��>
�.�|#��!�YPؾY���������|��wC���y�̽���S1�ZMݼ7���x   x   e����r��Rd��ZR�����2ܽb#�1�D�@�x�u;���v���9ɾ1�ܾ��=��:����1�ܾ�9ɾ�v��s;��C�x�4�D�h#�$ܽ����}ZR�od�hs��g���x   x   c2ݼ�\�vK=��j�� ���P���: � �K���z�9-���ɫ�쀿���ξ	�ؾz�۾
�ؾ��ξ耿��ɫ�=-����z���K��: ��P��& ���j��OK=�w\�2ݼ�qʼx   x   �:1��HR��e��̮��,ڽ:��:X0�YY��a��뗾M���4���Ⱦd6ξf6ξ�Ⱦ
4��O���뗾�a��YY�BX0�?��4ڽ�����e���HR��:1��Z!��Z!�x   x   e݉��暽�����ٽ�T�k�#��BG�b�n������П� m���B��Ⱦs!˾Ⱦ�B��!m���П�����c�n��BG�j�#��T���ٽ����暽U݉��g����z��g��x   x   ��̽��۽�?�����֜#��A���d�^ۅ�ȫ��-I���
���wǾ�x;�x;�wǾ�
��(I��ǫ��aۅ���d��A�ܜ#�����?����۽Ô̽��ý�(���(��m�ýx   x   ��E��. �P0��=G���d�n	���9��Wl��Qֻ��ɾ �Ҿ�վ�Ҿ�ɾSֻ�[l���9��g	����d��=G�P0��. �B���jL�8��s�<��pL�x   x   �`C��D��K��NY���n��م�9��@���d��"V̾�ؾ�M޾�M޾�ؾ!V̾�d��<��9���م���n��NY��K��D��`C�t�D��UG�LI�II��UG�w�D�x   x   ��|�f�x�n�z��[��>틾����k���d���m;Dg۾\��;��T��Eg۾�m;�d���k�����9틾�[��p�z�j�x��|����+��2	�����2	��'�����x   x   蜾�.��#���䗾_͟��G���ֻ��V̾ h۾��������쾺�� h۾�V̾�ֻ��G��_͟��䗾~#���.��蜾���,����#�����������#��*������x   x   击��h������ѯ���i��`
���ɾ�ؾ7��� ����� �2�侰ؾ�ɾ`
���i��ί�������h��ㇻ��MȾJ�վ��ྮ���n뾦�辿��L�վ�MȾx   x   �=ؾ+ɾ�v��.��W@��wxǾ�ҾQ޾d��R�O�f��"Q޾��ҾxxǾW@��.���v��+ɾ�=ؾ���TR������� ���������XR�����x   x   ��ٻܾ�ξ�Ⱦ�Ⱦ�z;��վvR޾͒�y��ђ�tR޾��վ�z;�Ⱦ�Ⱦ�ξۻܾ��O��-G���l�)��0�^�2� �0�l�)���.G�R��x   x   /�c��Rzؾ[2ξl!˾�{;	�Ҿ�ؾ�l۾�l۾ؾ�Ҿ�{;h!˾_2ξVzؾ^��.�����"�z�3�s�B��"N��(T��(T��"N�x�B�z�3��"����x   x   5%�����۾�3ξRȾ+|Ǿ��ɾ�\̾bt;�\̾��ɾ'|ǾRȾ�3ξ �۾���8%������/�//E��%Y��ri��$t���w��$t��ri��%Y�3/E���/����x   x   �6
�2��}ؾnȾ E�� ��%ݻ��k���k��'ݻ���!E��oȾ}ؾ5��6
�u��W�7�l�Q�:�j�79��gU����������hU��99��7�j�i�Q�W�7�w��x   x   �&�֬�P�ξ4���p��O���s�����s��O���p��4��M�ξլ��&�t��ʱ:��$X�1�u����������隿�o���隿��������5�u��$X�ȱ:�s��x   x   y���ܾ!~��{���K՟�7���&A��)A��:���I՟�w���%~����ܾy�w����7�L&X�̮y���������`W���ݪ��ݪ�cW����������̮y�N&X���7�v��x   x   ��D4ɾuȫ�F헾����ⅾ%��ⅾ����L헾vȫ�@4ɾ��S��n�/�o�Q�b�u�����H����ܪ�)���y���#����ܪ�J�������`�u�n�Q�o�/�S��x   x   (Iؾ@s��N-�� e����n�:�d�6�d���n��d��J-��Bs��+IؾI��S�"�z5E�L�j�Q��������ݪ������ռ��ռ������ݪ�����R���M�j�z5E�Q�"�J��x   x   i����9��[�z�T`Y��MG���A��MG�W`Y�\�z��9��f���|�꾵N���3�	.Y�l=�������Z�������ּ����ּ������Z������l=��	.Y���3��N�|��x   x   ������x��K�V`0���#���#�P`0��K���x�����\Ⱦ�b���~�B�e}i��Z����⪿J���Vؼ�Sؼ�H����⪿��Z��d}i�~�B���b��\Ⱦx   x   ��|���D�@ ���� `����@ ���D���|�߽��}�վz�c�)��.N�P1t�F���	v���㪿!���l���'����㪿v��G���P1t��.N�c�)�{���վڽ��x   x   �wC��&��\���ڽ�ڽ�\��y&��wC�r&��弬�S������0��6T�\�w�1����(^��s⪿o⪿&^���3���\�w��6T���0����O�漬�u&��x   x   ���7ܽ*-������.-��>ܽ���1�D��"��<6��X��`��-
3��7T�h4t�z]��}���������������~���x]��d4t��7T�0
3�b��W��<6���"��-�D�x   x   L�̽�����w���w������X�̽a�KpG����|Ѷ�-��,����0�a2N� �i�zA������9 ��: ������xA��%�i�d2N���0�+��&�뾁Ѷ����KpG�&a�x   x   t���lR��d=�HlR�m���	Ľɧ�!I��0��EҶ������!�)��B��5Y�;�j�{�u���y�v�u�?�j��5Y��B�!�)������HҶ��0��!I����Ľx   x   ]1��t�tt�]1����MI����r!I����o8��r��!���Z�3�I>E�,�Q��2X��2X�-�Q�F>E�[�3����!�n�j8�����z!I���WI�����x   x   ]ݼ���R]ݼ�z!���z��H�����AqG�$�����͝վ k��ET���"�k�/�?�7���:�?�7�i�/���"�FT��j��ϝվ	���	$��BqG�����H����z��z!�x   x   6ʐ�Gʐ���ʼ�w!�U}��}Ľ�`�/�D�,(��I���bȾ������C������������E��������bȾG���-(��'�D��`��ĽH}���w!���ʼx   x   � ��U������6:��ю��mҽ�>���G�c����柾5Ͼ���۾����F����	�����	�B��������۾1Ͼ��柾b�����G��>��mҽ�ю��6:����J���x   x   �顼�˼*���S�����\|ؽ�?���@��Xs��ݓ��_��Eoľ�d׾�����������侦d׾Foľ�_���ݓ��Xs���@��?�Z|ؽ������S�"*��˼�顼x   x   He�q!���;�4}��-����你:��W=���h��s��/^������r���4�Ⱦ��˾1�Ⱦy�������-^���s����h��W=��:����-��M}���;�a!��d<޼x   x   :���S�"}����uFŽ������b�>�H�d�����/��舤��ծ��6���6���ծ�判�/������J�d�d�>��������FŽe���(}���S�-:�[.�8.�x   x   輎�J���{!��@Ž�4�V��Y�'��G�h�%���b��Q���Zा�[��VाP����b��'��h��G�U�'�Q���4�@Ž�!��F���ڼ��?��yO��O��x   x   HOҽ�bؽ��m����& ��>9�V�U��s�f������TV��)�'�[V�����`����s�Y�U��>9�#& ���h�� �佄bؽJOҽL�Ͻ2HϽ-HϽ8�Ͻx   x   G*��-��,�b���'��;9���O���i��3�������������L�����|���!����3����i���O��;9��'�b���,��-�L*�|s�i��#W�q��~s�x   x   n�G�J�@�wE=���>��F�r�U�´i�y���㞌��\��l��K���O���l���\��㞌�u���´i�w�U�"�F��>�sE=�H�@�r�G���O��NV��%Z��%Z��NV���O�x   x   {뀾i=s��h�>|d�j�g��s�%2�������*���(��z.��L��r.���(���*������(2���s�_�g�;|d�߭h�n=s�z뀾�ˈ��������6���������ˈ�x   x   1ԟ�rΓ��g���L��&���ƌ���\��)��0,����
��3,��)���\��ǌ��"���N����g��sΓ�/ԟ�����ԝ��c�����ƾ��ƾg���ѝ������x   x   ܺ��	O��Q���%���\���������cl��B/�����qά����?/��cl����������\���%���P��
O��غ��ݝѾ���ѣ�����[������֣򾹯�ڝѾx   x   �۾{]ľ�����������S�����n����M��y��t���M��q�������S��£��������x]ľ�۾9��.I��p�`��t2�w2�a���p�0I�9��x   x   ;����R׾����̮�{ۤ���uM��]����0���.���0��\���rM����uۤ��̮�����R׾;�����
��Z���*�Yg7���?��|B���?�Xg7���*��Z���
�x   x   ��6��x�Ⱦ�.���W���򠾒��	o��Q,��P,��o��������W���.��}�Ⱦ0������� �,���@�Y�R�l�_���f���f�l�_�^�R���@��,����x   x   ��	�-���˾�/���ݤ��V������`���.���`������V���ݤ��/��
�˾.�뾼�	�3,!��A:��gS��vj�� }�^����ņ�`���� }��vj��gS��A:�1,!�x   x   ����� �ȾЮ�����h�������\���]�������f�������Ю��Ⱦ��뾛��
&���B�֤`�V>}�� ��W)��{	��z	��Y)��� ��Q>}�Ԥ`���B��
&�x   x   v�	����򰿾����Ob�������7�������7������Ob�����������s�	��&�g�E�^�g�����P
���{��u���*j��r����{��Q
������\�g�c�E��&�x   x   ]��zY׾�U,������#s��i��i��#s����P,��򏱾~Y׾_��4/!�/�B�֕g�*����͘�oo��C���������F���lo���͘�+���ڕg�1�B�2/!�x   x   ����YfľAY��l���$h���U���O���U�h�r���AY��Vfľ����E��:F:��`�M����Θ�0��2��o�ÿ[ǿi�ÿ4�� 0���Θ�L����`�<F:�G��x   x   H�۾GY���p���d��G�=G9�:G9��G��d��p��IY��H�۾��
���,��nS��D}�=���q��z���ƿ��Ϳ��Ϳ	�ƿw���q��>���D}��nS���,���
�x   x   tǾ�Wٓ�L�h�T�>�~�'��/ �v�'�X�>�P�h�Yٓ�tǾ�VG���b�A��j�k���������)�ÿ0�Ϳ�bѿ0�Ϳ)�ÿ�������l���j�A��b�UG��x   x   8៾Ss�W=�U��������R��W=�Ss�5៾$�Ѿ�Q�h�*� �R�,}�</��,����$���ǿ��Ϳ��Ϳ�ǿ�$��-���;/��,}��R�g�*��Q�$�Ѿx   x   ���y�@�B<�S���E�A��J<�y�@����ˬ����/{�s7�f�_�Q������-q��D&���ÿA�ƿ�ÿB&��)q�����R���i�_�s7�-{����ˬ�x   x   {�G��?����VSŽUSŽ��作?�|�G�fڈ�~������g���?��f�~͆����|����������������������}͆��f��?�j�����~���jڈ�x   x   >��ؽ�6������6���ؽ>�a�O��ҏ�-���E����?��B�b�f����:2��x���xw��,7��{w��x���82�����c�f���B��?�A���+����ҏ�]�O�x   x   FoҽL���=%}�+%}�E���Uoҽ*��EkV����� �ƾ� ��@�n�?���_��2}�
��(��֘�֘�'���	���2}���_�i�?��@�� �&�ƾ����DkV�6��x   x   >Վ�[�S���;��S�6Վ�pн����CZ�YI��2�ƾ��� ���w7���R�ڈj�)P}�$�������!���/P}�ڈj���R��w7�"�����3�ƾQI���CZ����oнx   x   �>:�B8�8��>:�S(���kϽo�}DZ����1�����S�]�*�#A��xS�u�`��g��g�v�`��xS�&A�]�*�S����+���!����DZ�o��kϽT(��x   x   +���˼Z��/.�^h��ekϽ:���mV�nՏ��������W�ui�^�,��P:���B�1�E���B��P:�^�,�ui� W��������pՏ��mV�*��mkϽ\h���..�x   x   ��������c޼j,.��&���н0����O��݈�[Ь��Ѿ%R��ư
����d9!�:&�7&�c9!����°
�)R���ѾXЬ��݈���O�9���н�&��},.�Rc޼x   x   ~?��%��<���E�8��p�ٽ$����L�I���\D���}¾ף߾����R�'��<�'�L�����ܣ߾�}¾]D��H�����L�"��Z�ٽ4����E��%��x   x   ;��f8޼_����X�9ؚ�zLؽ�r�ne?��q��L���_���¾k�Ծ���h��^�����n�Ծ�¾�_���L���q�he?��r��Lؽ=ؚ���X�g���8޼V��x   x   ]������>���y�Z���L�ڽy���3���\��(���薾����t��6罾Z���4罾�t������薾�(����\���3�|�?�ڽZ�����y���>���=������x   x   �gE���X�@�y�+6��7��������8�+�pNM��n����j���3������%���1���h�������n�vNM�<�+�������7��6��<�y���X��gE�7f<�#f<�x   x   /���!Ś������/���Gѽ����M�ħ)���D��D_��w���"����������󄾼w��D_���D�ħ)�M������Gѽ�/������*Ś�����P��㕑��P��x   x   �ٽ�/ؽ��ڽ3}�����b�a��|B-�*:C�'�X���j�~rx������rx���j� �X�0:C�yB-�_���b�+���*}㽼�ڽ�/ؽ߅ٽ�'ܽm
޽i
޽�'ܽx   x   ^w��^�t��-���E�����%��46�@H�j.Y��Kg��p���s��p��Kg�r.Y�>H��46���%����E�*��z���^�_w�v�!�"��Y$�+�"�v�x   x   o�L�L?�֟3�z�+���)�.<-�J26���B�*YQ�v�^�Xgi�o�o�\gi�~�^�+YQ���B�F26�/<-��)���+�֟3�L?�w�L���Y���c��zi��zi���c���Y�x   x   �僾��p���\�J;M� �D��1C��H��WQ��x\���f�E�m�c�p�?�m���f��x\��WQ��H��1C��D�E;M���\��p��僾���`��K�������K����`����x   x   �/��q;��8��*�n��5_��{X�G)Y�X�^�O�f�v�m��r��r�t�m�Q�f�d�^�E)Y��{X��5_�-�n�:��r;���/�����þ�:ξ�0Ծ�0Ծ�:ξ�þ��x   x   >g¾=L��hٖ�]����w��j��Fg�{ei�$�m��r��s��r�#�m�{ei��Fg��j��w�\���gٖ�@L��8g¾�ھU�ﾪ� �	��5������ �R���ھx   x   ��߾.������dx���넾�hx���p�o�)�p��r��r�*�p�o���p�ix��넾fx�����'�����߾A����@�@'�Y�$���)���)�X�$�>'��@�=���x   x   ������Ծid��\���n��������s�Lo�9�m���m�>�m�Ko���s����f���X���ed����Ծ��������#���4���B��L�j9O��L���B���4��#����x   x   � �&��Y׽�灡������4�p��hi��f��f��hi�0�p����������b׽�!�ᾡ ��?��%5�*�K�Et_���m���u���u���m�Lt_�%�K��%5��?�x   x   �����y����������omx�wKg���^�*}\���^��Kg�omx����􂡾i�����辴�1�&��(C��*_�=�x���7�������7��썆�=�x��*_��(C�,�&�x   x   (1��辻ٽ�R���*��j��/Y��]Q��]Q��/Y���j�*P����ٽ���(1���+�wL��m��3��P�������������������Q����3���m�L���+�x   x   r�f��i��}���w���X�SH���B�ZH���X��w�}���h��^��o���+��O��It������F������ᄳ����ބ�������F�������It��O���+�x   x   ��A�Ծ-��V���^@_��:C��96��96��:C�]@_�R���1��F�Ծ��E�&��L�Kt������P���/��L����:ƿ�:ƿP����/���P������$Kt�L�B�&�x   x   �������7ᖾ��n�q�D�$E-���%�)E-�n�D���n�4ᖾ��������D�f-C�nm�o����Q��*��ƿ�`п��ӿ�`пƿ/���Q��m���lm�e-C��D�x   x   �߾MV���"��^IM��)��������)�SIM��"��QV���߾���a,5��1_�U7���I��,2��_ƿ��ӿOBۿQBۿ��ӿ\ƿ+2���I��U7���1_�`,5����x   x   �s¾*F��	�\��+��O�Ki��O��+��\�*F���s¾����#�"�K���x� ���Ū�:����cп�Cۿi	߿�Cۿ�cп:���Ū� �����x�"�K��#����x   x   &=��Uq�b�3�c������ġ��a��`�3�Tq�#=��!ھ�I��4��_����ճ������\@ƿ'�ӿoEۿlEۿ%�ӿ`@ƿ����ҳ������_��4��I�}!ھx   x   u��_?�7�ّ�WTѽő�:��_?�x��.��*�,2�E�B�h�m�?��[ �������Aƿ�fпo�ӿ�fп�Aƿ����] ��?��k�m�H�B�(2�*��.��x   x   ��L�@p�k�ڽ@��@��z�ڽAp���L���j%þ�� ��$�!L���u�w���{��t���J����ƿ�ƿG���y���}��u���~�u�L�	�$��� �l%þ��x   x   |���Lؽ!���4B��'���zLؽ~����Y��q���OξW��&�)�\IO��u��@������ɪ�`8���"��d8���ɪ�����@���u�dIO�&�)�U���Oξ�q����Y�x   x   Y�ٽ�ۚ�]�y�K�y��ۚ�l�ٽ����	d����LGԾ���<�)��L��m��������2P���Y���Y��2P����������m��L�8�)����RGԾ���	d����x   x   ���8Y���>�GY����OKܽ��"�Ԛi��Ѡ��HԾ����$�;�B�ކ_��x��=��ᓌ�Î�ݓ���=���x�ֆ_�?�B�"�$�����HԾ�Ѡ�Ӛi���"�UKܽx   x   ��E���������E��j���/޽As$���i�ߦ��YSξ�� ��6���4��K�=_�m��Zt��Zt�m�=_��K���4��6��� �SSξ榞��i�Hs$��/޽�j��x   x   �[Q޼�@�<�[���N0޽��"��d�"u���*þ�
��O��&#�=65�G9C��L��(O��L�J9C�=65��&#��O��
��*þ!u���d���"�P0޽b���5�<�x   x   -��>-������Z�<�)j��NLܽݎ���Y�i���5��%+ھ̼��!���N���&��+� �+���&��N���м��)+ھ�5��i����Y���eLܽj��c�<�����x   x   Bn��rYͼ9�Q��.��;t�h��HQ�Mf���꥾
Ož\�⾮���������7������������e��Ož�꥾Mf���HQ�h� tེ.��Q�9�vYͼx   x   4Lͼ���k� �u�_����jٽ�h�z�>���o�M�����X����Ҿ�߾t�tt��߾��ҾX�����M���o�r�>��h�3jٽ�����_�`� ����nLͼx   x   i(��� �}�C���y�����a}Խ�	���,��T��{�QҐ��I������%��g긾�%������I��UҐ�"�{��T���,��	�Y}Խ������y�v�C��� �N(����x   x   o�P��_�X�y�xא�཭�fԽE�^3��f<���Z���v��&�����������������&����v���Z��f<�d3�E�fԽ߽���א�C�y���_���P��IJ��IJ�x   x   1��l������뵭�AQ���_۽j���a*�0�*�	WA�\�U���e��6p�n�s��6p���e�S�U�	WA�4�*�`*�d���q_۽LQ��絭�����������˚��ښ��˚�x   x   ZP�Kٽ�dԽ>UԽW۽�꽸� ����.
 �cb0�5�>��bI�oO�oO��bI�2�>�eb0�5
 ������ �'��W۽3UԽ�dԽKٽVP�������꽾��x   x   �O��S�I	��7������� ����J�@��7;'�1��7���9��7��1�A;'�6��J������ ������7�S	��S��O�k!%��)+��M-��)+�_!%�x   x   �)Q��>�A�,��!� �2���F�V!��h�X%$��~*��.��.��~*�\%$��h�`!��F�/��%��!�B�,��>��)Q���a�în���u���u�ˮn���a�x   x   mS���o�Q�S�Q<���*�   �����f��( ��$��f(���)��f(��$��( ��f����"  ���*�wQ<�E�S��o�pS��x듾����E��J̨��E�����|듾x   x   �ԥ�	:����{��Z�EA��V0�=4'��!$���$�c�&�bK(�gK(�\�&���$��!$�=4'��V0�EA��Z���{�	:���ԥ�������ʾ_�׾Z޾Z޾]�׾��ʾ����x   x   �6ž�������v��U�]�>�w1�8{*�Ee(� K(�{v(�!K(�Ie(�7{*�q1�U�>��U���v�����񩾵6ž�_�  ��[Z�!�������eZ� ���_�x   x   <z⾳A��a7�������e��UI�z�7�Y	.���)�K(�{K(���)�U	.�y�7�VI���e����`7���A��Az�����T�Ry!���+�hJ1�kJ1���+�Ny!��T����x   x   |�����Ҿ%�������V#p�O���9�
.�\f(�0�&�af(�
.��9�O�L#p����������Ҿ���wt�p�(�^�;� �J���T��DX���T���J�^�;�n�(�xt�x   x   ���2�߾���.�����s�GO�f�7�^}*���$���$�Z}*�_�7�CO���s�5������/�߾���.'!��;��S��h���w�Q��F����w�$�h��S��;�1'!�x   x   =��i^�&ٸ�'���>&p�xYI��	1�%$��* �%$��	1�|YI�B&p�$���ٸ�e^�>��-�*��pI�efg�T;��6��(�� ���-��2��T;��nfg��pI�&�*�x   x   w���_����P���H�e���>��8'��i��i��8'���>�C�e�L������_�z��,�/���R��u�m��Ŭ��'��:���:���'��Ƭ��m���u���R�/�/�x   x   ���d�߾��������U�]0����$����]0���U������\�߾���>�/�N�U��}�������������׺�c���׺�������������}�D�U�A�/�x   x   K��F�Ҿ�=����v�0NA� �YK�VK� �,NA���v��=��K�ҾO��N�*�;�R�%}��4������ea���[ǿT?οZ?ο�[ǿ_a�������4��+}�@�R�J�*�x   x   ���?J���Ȑ�1�Z�C�*�Ř����Ș�C�*�B�Z�~Ȑ�>J�����!,!��uI���u�a���¾��
e��|�Ϳ0�ؿf{ܿ(�ؿ~�Ϳe������_�����u��uI�&,!�x   x   Å⾵�����{�J^<�L'�P� �K� �R'�<^<���{���������z��$;��mg��p��(����c����Ϳ�bܿ�俱��bܿ��Ϳ�c��+����p���mg��$;��z�x   x   ~Cž�D����S�!.�����3�꽶���'.���S��D��~Cžl��Ԯ(�I�S�;@������į���_ǿ1�ؿH俻��H�1�ؿ�_ǿů������;@��H�S�Ԯ(�l��x   x   2⥾��o��,��B�d۽ d۽�B��,���o�0⥾�o��]���;�ӎh���y-���ݺ� Eο�ܿ�	��	��ܿEο�ݺ�u-����Ҏh���;��]��o�x   x   R`����>�N	�fgԽ�Z��YgԽR	���>�V`���ι�o����!��	K�'�w��%�����!��}Fο>�ؿ�gܿF�ؿ{Fο�� ����%��)�w��	K���!�k���ι�x   x   BAQ��d�|Խ�í��í�+|Խ�d�FAQ������˾�e��+�[�T�`���L����຿dǿ�ο�οdǿ�຿O���엕�]��W�T��+��e��˾����x   x   d��gٽ桢��ᐽ롢�cgٽd�Nb�l���׾���Y1�~UX�8���'���0������[j���l��`j�������0���'��;���UX�Y1����߶׾f��Tb�x   x   !q�[!���y��y�n!��7qད8%���n�eY���q޾���EZ1�5�T�"�w�I������唣��ƨ��ƨ�唣�����L��&�w�)�T�AZ1�����q޾pY����n��8%�x   x   /����_���C���_��.��a��C+��u�-ᨾ/s޾���a�+�K���h�fE��'w��7����=��3���*w��fE����h�"K�h�+����+s޾ᨾ�u�C+�m��x   x   eQ��� ��� �yQ��暽'�꽬h-�p�u�z[���׾ i���!�6�;��S��yg��u��)}��)}���u��yg��S�6�;���!�i���׾�[��|�u��h-��꽉暽x   x   T>����/>��mJ�~�������D+���n�S��!˾���qd�Y�(��/;���I���R�~�U��R���I��/;�Z�(�od����,˾O����n��D+���꽏����mJ�x   x   &aͼ\aͼ[��mlJ��暽��潷;%��b� ���ֹ��zྡྷ����7!���*�J0�I0���*�7!�������z�~ֹ�
 ���b��;%���潎暽hlJ�S��x   x   n�ȼԧ��$���Z��埽D����^�S�ju���ᦾ�%ƾ�G�b\�����&��� �+�����i\���G�y%ƾ�ᦾku��j�S���(��埽��Z�%�ާ�x   x   i�����5�(� �e������ٽO��fx=�&�m�mϏ��������о?�ܾ����E�ܾ�о������nϏ�0�m�^x=�I���ٽ���7�e��(�������x   x   ����(���H��\z�����b�Ͻ�(�Kh'���L��s�����󐛾Tݧ�����Q�����Uݧ�������s���L�Eh'� )�a�Ͻᐠ��\z���H��(���w�x   x   �Z���e��Nz��捽 ঽ<ɽK������y/�A~K�t�e��X{�㇅�"���+���݇���X{���e�/~K�y/����S���4ɽ�ߦ��捽�Nz���e��Z�ӼU��U�x   x   {̟��垽O����צ�᳽��Ƚ=g�=5�����+���<�PK�Z6T��_W�P6T�cK���<��+����:5�/g彀�Ƚ&᳽�צ�D����垽^̟��>��㡽�>��x   x   ��佄�ٽ��Ͻnɽ��Ƚ��Ͻ��޽��"<�=��ng���&���+���+���&�lg�A��&<�ۥ���޽��Ͻ��Ƚ`ɽ��Ͻ��ٽ���d;v�v�[;�x   x   ���������f��7U�e�޽�]�h<�i��������	��F�����F���	���W���`<��]�Y�޽)U当f����������4l)���0�
53���0�"l)�x   x   �dS��[=�ZP'����(����25��署�����������������������5��/5齯��(���YP'��[=�eS���f��Yu��}��}��Yu���f�x   x   �a��z|m�ܺL�b/�ń��0�����s��Z��꽶,��,��Y��m�뽐����0�̄�b/�кL��|m��a������9좾�䪾�����䪾8좾����x   x   �ʦ�t���/�r��cK��+�������S���4��'��4��&����^�������+��cK�:�r�r����ʦ����bϾy
ݾs@侁@�s
ݾbϾ���x   x   6ƾ������She�]�<��X�r�	�l���(콾���5����)(�h���m�	��X�T�<�Zhe�������.ƾuz�����h	��&�{��&�h	�����jz�x   x   �,����y}��:{���J�O�&�R=�&���M��彥��@����T=�W�&���J�(:{�w}�������,�>^�R��7�$�k�/�-_5�._5�f�/�2�$�Y��>^�x   x   @����Ͼqɧ�nx���T�n�+�`�������(�t���(�����f��i�+��T�fx��hɧ���Ͼ@�����b+�S?�J,O�1eY���\�;eY�H,O�S?��b+���x   x   r����ܾ]������XJW�g�+��>������꽴������>�c�+�^JW����l�����ܾm����"��=�
[W�)�l���|�;���4�����|�0�l�[W� �=���"�x   x   ���k㾹>������n"T��&�؝	�k�/��s�ߝ	�%�&�r"T�󕉾�>���k�����,��UL�LKk�����T����╿�a���╿Q�������VKk��UL���,�x   x   O���l㾒����z����J��\������������\���J��z�������l�S���1�yvU���y��Ӎ��a�����z���z�������a���Ӎ���y��vU��1�x   x   ����ܾ�ͧ�	B{��<����������罺�������<�B{��ͧ��ܾ�����1���X���� e���O��Ҫ�����34�����ժ���O��#e������X���1�x   x   ���- оg����re��+�M6�:�:�K6��+�yre�h���4 о���ő,�yU�䎀�����h���m����ʿS�ѿZ�ѿ��ʿ	m��e�������玀�yU�,�x   x   hI��i���F���oK�
��f��(`�j����oK�D���j���aI����"��ZL���y��f������+t��i7ѿkܿ&�߿cܿk7ѿ4t�������f����y��ZL���"�x   x   8�B���s��m/��/���޽�޽�/��m/��s�E��8����=��Rk�t׍�S���o���8ѿ��߿�p��p習�߿�8ѿ�o��S��s׍��Rk��=���x   x   �ƾ�ŏ���L�5���b彈�Ͻ�b�8����L��ŏ��ƾ�e��j+�RdW������f������̔ʿpܿxr��`�xr�pܿ̔ʿ�����f������QdW��j+��e�x   x   ئ�1�m�k_'�xz����Ƚ��Ƚdz��p_'�7�m�ئ�z�㾯���]?��m�����A��e ���ѿ��߿t�t���߿�ѿg ��<�������m��]?����w��x   x   �n���n=��#��ɽ*賽�ɽ�#��n=��n��C���m�����$�49O���|��ꕿn��� <����ѿ�ܿK�߿�ܿ��ѿ�;��q����ꕿ��|�99O���$�f���E���x   x   �|S������Ͻ�㦽�㦽��Ͻ����|S����-uϾ|s	���/�9tY������j������
���ʿ�>ѿ�>ѿ�ʿ�������j������4tY���/��s	�1uϾ���x   x   ޮ�e�ٽ`����g���D�ٽޮ�1�f����P ݾ�3�n5���\�g����앿�������v��1|��$v����������앿j�����\�n5��3�F ݾ ���<�f�x   x   ������gz�hgz�0����彚�)�yu������X�2��Ko5�.wY��|�����Ql���Y�����������Y��Ql�������|� wY�Go5�6���X侏���yu���)�x   x   T埽��e�R�H�~�e�:埽m`�0��:}����Z侤5�*�/��>O��m�ؚ�� ލ��n��ѱ���n��#ލ�ؚ���m��>O�3�/��5�Z������:}���0�}`�x   x   ֮Z�>�(�n�(��Z��Y�����|P3�h<}������$ݾ/w	� �$�Ce?�@nW�_k�g�y�V���\���l�y��^k�EnW�Ce?���$�)w	��$ݾ����v<}��P3�u���Y��x   x   �)�+���)�^�U�h�������0��}u�T�� |Ͼl�������s+�.>��gL�I�U�6�X�?�U��gL�0>��s+����m���|ϾN���}u���0�������d�U�x   x   @�ἀ��Ջ���U�NZ���c�e�)�p�f�⸖��ȼ�?��`m��&�E�"��,���1���1��,�I�"�~&�am�H���ȼ�޸��w�f�w�)��c�EZ��r�U����x   x   �6ټ�|��X��`����>�՗�͗R�ކ���q���1ľ!�ྷ{���9�4�?�$4��9��{��.�ྑ1ľ�q��߆��ؗR�ȗ��>�����`�Y��|�x   x   4o�d�	�_.�A9i��1���Wؽ���k:��Ni�0��Ĵ�������˾�%ؾY�޾N�޾�%ؾ��˾���Ĵ��2���Ni��k:����Wؽ�1��Z9i��^.�<�	�zo�x   x   �G��T.��K�z�y���xʽ��ɸ!��E��'j��������ύ���
��_����
��ҍ����������'j�ՁE���!���xʽ��q�y��K��T.��G�o3�x   x   �`� i�`�y�T���砽͒��r���
���$�b�>���V��Qk��
z�4���?����
z��Qk���V�P�>���$�	�
�{�Ò���砽r��?�y�~ i�/�`��!]�""]�x   x   T�����4����ޠ�Gש������ѽ��ｬ��G���)�2M6��>�rWA��>�FM6�Ӡ)�A��������}�ѽ���\ש��ޠ�$�����7��]�������O���x   x   潻6ؽ�]ʽ����y��ԓ��DĽӽV�F��[f��r��?��?��r�]f�F��]��ӽDĽ񓻽}�������]ʽ�6ؽ���1��V���V���1�x   x   )~�2��������ѽ;Ľ�侽���פǽ2ѽ�ڽo��=�⽇���ڽBѽΤǽ���徽;Ľ�ѽ����1��~���*���2�wV5���2���*�x   x   �vR��N:�T�!���
�3��ӽp����O��t������Ɛ��xk��`k��ϐ�����g����O��n���ӽ<����
�R�!��N:�wR��g��
w�qM�ZM�w��g�x   x   �r��T+i�dE��y$�������ǽ����tp��:����z��s3���z��>���pp�������ǽ������y$�dE�e+i�s������w����﫾�Ү��﫾x�������x   x   �Z���Ij�ނ>����L)�� �н^쵽t𥽤����+���+������m�l쵽(�нc)�����ڂ>�Uj���Z���M����Ͼ��ݾ'V�4V���ݾ��Ͼ�M��x   x   �ľ@���p��V�V��)�MV�.ڽՄ��u���)���
���)��3u��Є��"ڽBV���)�a�V�p��A����ľ���[����	������������	�T���x��x   x   ���� ��q��� 2k�-56��a��~��^���,��8)��-)���,���^���~��a�956�2k�m���� �����:�����R�$���/���5���5���/�M�$���:��x   x   �^��͑˾9y��|�y��h>�/����_���t��G����t�� _�����/��h>�n�y�3y��ݑ˾�^��5���*��
?��O�#GY��\�-GY��O��
?���*�5�x   x   0+��ؾ����AЀ�@A��/����煸�c諒X諒څ������/�@A�GЀ������ؾ*+���!��/=���V�jl�5|�JF��CF��5|�jl���V��/=���!�x   x   �%�*�޾����р�5k>�'d�pڽb��m��f��ڽ2d�5k>�р�����%�޾�%��T+�4^K�6dj�'���$��TK���ė�ZK���$��'��@dj�/^K��T+�x   x   n1�~�޾����0�y��96��Y�5�н��������-�н�Y��96�.�y�������޾q1��R0��[T�{x�B+��2����)�����������)��2���?+�� {x��[T��R0�x   x   �'��ؾQ}��f9k��)��1����ǽuM����ǽ�1���)�v9k�H}���ؾ�'��S0�$qW�f��杓��U��)��ƪ���׿�����,���U��靓�`��qW��S0�x   x   i.�-�˾#�����V������c���j����彌����V�#���5�˾n.��W+�^T�����֕��s��=��k�ȿ��Ͽ��Ͽn�ȿ5���s���֕����^T��W+�x   x   1h������v��q�>�X��5ӽ^侽:ӽR���>��v�����*h��u�!�cK��x�����u������zϿ�"ڿ��ݿ�"ڿ�zϿ���t�������x�cK�{�!�x   x   ���ħ��oj�ބ$���� @Ľ@Ľ���؄$�mj�ŧ�����Y;��6=�Wkj��.���X�����<|Ͽ��ݿ)<�,<忯�ݿ6|Ͽ����X���.��Zkj��6=�R;�x   x   x$ľ����SsE�2�
�+�ѽ���-�ѽ2�
�QsE�����{$ľ�����*���V������΃��h�ȿ�%ڿ�=�鿼=��%ڿh�ȿ΃���������V���*����x   x   �g���?i���!�;��������*�潺�!��?i��g��W��?���?��ul�:+���/������Y�Ͽh�ݿY?�V?�d�ݿ^�Ͽ�����/��;+���ul��?�D��V��x   x   ���za:���9����ܩ�2�����ha:�����]��������$��O�)C|��R���ȫ��߿���Ͽ�(ڿN�ݿ�(ڿ��Ͽ�߿��ȫ��R��*C|��O���$������]��x   x   >�R����rʽ�頽�頽�rʽ��H�R�㴖���ϾG�	��/��UY�|N���͗��ɫ������ɿ��Ͽ��Ͽ�ɿ�����ɫ��͗�yN���UY��/�N�	���Ͼ㴖�x   x   ���Qؽ<�����C���Qؽ����g�,�����ݾe����5���\�XO���T��\3��ň��!�����&����Y3���T��[O����\���5�`����ݾ&�����g�x   x   E9潳0����y�o�y��0��X9��*�+*w�U��&n�����5��XY�DH|�/��h����_��}��}���_��g���/��IH|��XY���5���-n�d��$*w��*�x   x   ���X>i���K�?>i�����V�]�2��o�设�o�W����/�EO��}l�K��a5�������ߕ�����d5��J���}l�KO���/�W���o�设xo�_�2��V�x   x   U�`�.h.�]h.�q�`�xĤ��~���q5�-q�����ݾ�	��$�(?���V��wj�P�x�������U�x��wj���V�'?��$�
�	��ݾ���:q�r5��~��gĤ�x   x   X]�:
�]�XF]�ѥ������2�D/w�������Ͼ����G���*��A=�`pK�NmT�ЁW�EmT�`pK� B=��*�E��������Ͼ����4/w���2����$ѥ�`F]�x   x   ������H��E]�@Ť�qZ�!�*�L�g�����f�����v��E��!�	e+��b0��b0�e+��!�E�w������f�����V�g�0�*��Z�<Ť��E]��G�x   x   6x㼤�����!���a�K����⽠����M��=��I0��������ھ��Uy��A��;
��A�Ky�"�򾦹ھ����I0���=����M�������A����a���!�����x   x   �������e0�.~h�f蜽2�ӽ0�G�4��a�
_���/��̳�	�ľ��оs׾i׾��о�ľ̳��/��_��(�a�G�4�0�I�ӽj蜽J~h��e0�������x   x   �!�c[0�UYK��v�Q���Q�ý
��]��w�<�R�_��k��9�5���[���Σ��[���5��5�k��`�_�g�<�T����S�ýC����v�>YK�s[0��!�2�x   x   X�a��eh�� v��/��g������Uڽ�}�S8�>i2�pI��\�R�i�q�'q�K�i��\��I�-i2�P8��}�`ڽ���c���0��� v��eh�m�a�O]_�c]_�x   x   �����Ҝ��晽�x��݇���Z���#��M�ڽ�z���������	%��q,�u/��q,��	%��������z��J�ڽ�#���Z��ꇠ��x���晽Ӝ������e��ᯥ��e��x   x   x�⽱qӽS�ý���|Q��$���<j��Iҹ��eȽ��ؽ��罂��X��R�������罡�ؽ�eȽ5ҹ�Aj��G����Q�����^�ý�qӽu��7��������*��x   x   Or�������"�ٽ\��Ja��k��|��tڤ��5���)������1P������\)���5��oڤ�z|��/k��:a��@��"�ٽ������Er�~(�_i0�nO3�li0�q(�x   x   ��M�w�4����j���ڽ/����t��U���ƌ�B'���ꉽ�G���G��뉽Y'���ƌ�]���t��&�����ڽ�j���g�4���M�ec��Os�ͽ{���{��Os�
ec�x   x   <*��/�a�ܶ<�� �EW���MȽa̤�����m�{�T�k�H�c���a�T�c�W�k�@�{�����Z̤��MȽPW��� �˶<�>�a�=*�����򿠾�.�����.��񿠾���x   x   ����J���_��M2��m�?�ؽ
#����%�k�9�T��TJ��TJ��T�+�k���#��O�ؽ�m��M2�%�_��J������B����˾�پ,g�7g�	�پy�˾�B��x   x   qιt���X����H�~��������(މ�G�c��OJ��QB��OJ�b�c�%މ�������w�� �H��X��t��iιȄݾ����������4������������ݾx   x   `�ھ;���ڎ�t�[��$����|���:��p�a��MJ��MJ�g�a��9��}������#�$�u�[�ڎ�4���h�ھf� ��q��j!��=,� �1�!�1��=,��j!�r�e� �x   x   �z�X�ľ!��h�i��X,�C���+9��:��l�c�n�T�{�c�:��B9��2����X,�_�i�	!��e�ľ�z�I����&�o�:��oJ��xT�|�W��xT��oJ�n�:���&�K��x   x   �j���оWG����p�G�.�����푴�Mމ�r�k�u�k�Dމ�֑������W�.���p�bG���о�j�-��/�8���Q�}�f�J&v�y=~�m=~�E&v���f���Q�/�8�.��x   x   �3�U�־ۺ��A q��Z,�����������{����������Z,�5 q�ͺ��R�־�3���&�MgF��d�����{�� b���ē�b���{������d�IgF���&�x   x   C.
���־[I����i�&�$���罗%�����������%��w��"�$���i�iI����־E.
���+�
O��0r�w��9^������䦿䦿����9^��w���0r�O���+�x   x   o5�խо�$��]\���� �ؽ"Τ����!Τ��ؽ��i\��$��˭оl5���+��R�$Gy�ܤ�������?������z���?������ߤ��Gy��R���+�x   x   n�|�ľ�ߎ���H��s�uTȽ�t���t��kTȽ�s���H��ߎ���ľn��'��O��Hy��ő�����Gj��N�¿�Eɿ�EɿQ�¿Aj�������ő��Hy��O��'�x   x   ��� ���_���W2�d��vƹ��h���ƹ�d���W2��_��!��������lF�!5r����������;��k�ȿ�ӿ>�ֿ�ӿm�ȿ�;���������� 5r�lF���x   x   O�ھ�"����_��*���ڽ|d��gd����ڽ�*���_��"��K�ھk��Ѻ8��d�oz�������l����ȿ-uֿӜݿ՜ݿ1uֿ��ȿ�l������oz���d�Һ8�f��x   x   ���T��K�<�=t�����������:t�J�<��T������ ��'�]�Q����b��=D���¿�ӿQ�ݿ{C�Q�ݿ�ӿ�¿=D���b����^�Q��'��� �x   x   %&����a������ٽBX��TX����ٽ�����a�"&��'�ݾ�z���:���f��������f��&Kɿ��ֿٟݿ֟ݿ��ֿ+Kɿg�����������f���:��z�'�ݾx   x   }6��|�4������̋�������k�4��6��SR��q����u!�=|J��3v�Di��{릿\���Lɿ�ӿ�yֿ�ӿ�LɿT��}릿Fi���3v�A|J��u!�i���SR��x   x   �M�Y)��ý��������
�ý_)��M�峓��˾���J,��T�>M~�@͓��즿����¿8�ȿ2�ȿ�¿����즿=͓�8M~��T��J,����˾賓�x   x   �����ӽ����z6������x�ӽ����c�7Ѡ�Aھ_��x�1���W��N~�Bk��W����H���r��<C���r���H��T���?k���N~���W�v�1�[��8ھ/Ѡ��c�x   x   ����朽7v�+v��朽���/(� ns�5B���~�KB���1�։T��8v�U���h�����`���a������h��X����8v�ɉT���1�OB��~�DB���ms�/(�x   x   ���A�h��gK�1�h�{��ｖ�0�%�{��,��;��M��N,���J�r�f�$��Ԁ��?���AΑ�9���ր��$��i�f���J�"N,�N��6���,���{���0��x   x   u�a� n0�n0���a�N�������`j3���{��D���ھT�{!��:��Q��d�nCr��Xy��Xy�qCr��d��Q��:�{!�P��ھ�D����{�ij3�����B���x   x   ��!�u����!���_��˥�#����0�5ss��ՠ��˾��������'���8�yF�\%O��R�U%O� yF���8��'�������)�˾�ՠ�'ss���0�����˥�Ā_�x   x   \�������U1�]�_�N���ｃ3(���c�0���c[��T�ݾ^� ���V���'�J�+�G�+��'�[����_� �^�ݾ\[��-���c��3(��K���M�_�J1�x   x   `漁���� ���]������ڽ	c��.E�f{�v��la����о���i����$����Y����羫�оea��v��`{��.E�c���ڽ�����]��� �����x   x   �������>.���b�y����˽k���O,�8�V�����F��ت���\ƾEK̾=K̾\ƾت��F�����E�V��O,�h���˽x�����b��>.����V���x   x   �� ��4.�t�F��Pn�����e��2��b�D 2�t�R�h�q�ߩ���L�����r[������L��ک��g�q���R�7 2��b�2뽲e������Pn�:�F��4.��� �ة�x   x   а]�e�b��Cn�)����Β�}����̽�V�r�M�%���:�:]L��*Y�
�_�"�_��*Y�1]L��:�@�%�r��V��̽~���~Β�)����Cn���b��]���[���[�x   x   �l��圗�����\ƒ�@ʖ���������#�ǽ� ⽖(��J9�9|�I+��|�:+�C|�D9��(��� �'�ǽ��������Hʖ�^ƒ�믓�򜗽�l��R2������P2��x   x   ��ڽ��ʽ�L����������4��I�����:��sn��<ʽwԽ�oٽ�oٽ�ԽBʽqn���:���Q����4������	����L����ʽ��ڽ�1�N��Y���1�x   x   �J����?�x̽���������������c������P���V���Z䔽f���)��������c�����������������̽B�����J�(�!�68*��-�@8*�$�!�x   x   wE�4,��K��1�v�ǽ+ޤ����f�s�'e_�{%U�Q�P��O��O�\�P��%U�-e_�a�s����'ޤ���ǽ�1�K�4,��E�6uZ��(j��vr��vr��(j�7uZ�x   x   ��z���V��2�[���#���U��,Y_���<�: (�gv��D�ev�9 (�R�<�8Y_��U��#����[��2���V���z�����t��������������s������x   x   �뙾����F�R�x�%������Q���⌽�U���'�?h��A��A�4h���'�U��⌽�Q������q�%�U�R������뙾a�����þ�aѾ��ؾ��ؾ�aѾ�þb���x   x   I��Y1����q�A�:��"���ɽ����9�P��h��<�����<��h�:�P�������ɽ�"�M�:���q�X1���H���Ծ�p��>)��n
�9)�����pԾx   x   _�о����O����=L�d���ӽ���F�O��4�n:�_:��4�5�O������ӽ"d��=L�L�������e�о�+��aM����6%��*��*�4%����gM��+��x   x   1q�ֺ��8��>
Y����Lٽ�̔���O�'f�]`� f��O��̔��Lٽ��9
Y��8��ֺ�2q羼Q
������2��A�IK���N�IK��A���2�����Q
�x   x   ����Dƾ����'�_��d��Mٽ���N�P���'���'�C�P�����Mٽe�6�_�����Dƾ�������5�0��{H��\�1k��r���r�-k�%�\��{H�4�0����x   x   3���3̾H����_����ӽ����TU��<�CU����.�ӽ����_�H���3̾6�������=��WZ���s�����s��;���s��������s��WZ���=����x   x   ��5̾����ZY��g�r ʽp䌽S_�%S_�l䌽Z ʽ�g�[Y�����5̾��Q1$���E��g������������,���+���������������g���E�U1$�x   x   ����Gƾ:<��DL�_'�W��xV��=�s�zV��'W��_'�DL�3<���Gƾ���I2$�_�H���m�	���ׯ��X�������U������X��گ�������m�W�H�I2$�x   x   �����ۺ�m�����:��
��W(��������I(���
��{�:�o����ۺ���������E��m�@����<���쬿�_��bl��hl���_���쬿�<��B����m��E����x   x   �y�zȪ��q���%�q��⤽��#⤽g�ὖ�%��q�yȪ��y���%�=�g����=�������{ǿ��ʿ{ǿ������=����	g�#�=� ��x   x   ��о
:��ҶR�hd���ǽ����l�����ǽgd�ѶR�
:����о�W
�~�0�#^Z�	��������:����ʿ�7ѿ�7ѿ��ʿ6�������
���$^Z��0��W
�x   x   �T��ՙ��'2�@C�؟��24��ݟ��8C�%2�ՙ���T��99�����G�H�d�s���'\��%c���}ǿ�8ѿ��Կ�8ѿ�}ǿ%c��(\����d�s�G�H����89��x   x   ������V�AX��̽^���o����̽IX���V�����h+Ծ�U�y�2���\�O����������Jq����ʿO:ѿL:ѿ�ʿNq���������P�����\�x�2��U�j+Ծx   x   ��z�E,��$����1͖�����$�E,���z�:�����������A��k��y�����\\���r��I�ǿ�ʿP�ǿ�r��V\������y���k���A�������7���x   x   �$E�����^��ϒ�ϒ�_������$E�Ȫ����þ��S&%��VK�Һr����+���m����f��O��J���f��r���/������ͺr��VK�U&%�����þΪ��x   x   ]��˽꽓�Ը��⽓��˽]���Z������uѾ/5���*���N�h�r��{�������`��������������`�������{��l�r�ƢN���*�,5��uѾ|�����Z�x   x   ��ڽ�����Wn��Wn�������ڽ�"�Fj�Ǣ��ؾ�{
�Λ*�dYK��k�� ����������D���D���������� ���k�[YK�˛*��{
��ؾǢ�Fj��"�x   x   ���6�b�YG�2�b�	���T�NP*�ܖr� ����ؾ7��)%���A��\�	�s����Ɉ�ZƊ��Ɉ���
�s���\���A��)%�7���ؾ����זr�IP*�T�x   x   ;�]�RF.�NF.�V�]�zK����}4-���r�^ɢ�EzѾ���8����2���H��iZ��,g�g�m�p�m��,g��iZ���H���2�9�����@zѾiɢ���r��4-���uK��x   x   �� �S��k� ��\�"���	R*�#Kj�������þq�\�����0���=�5�E�ϴH�1�E���=���0����\�p��þ􈚾Kj��R*��%���|\�x   x   ���������!\��L��X�#"���Z��������?7ԾaH���`
�����*@$�&@$������`
�cH��G7Ծ���������Z�+"�5X罘L��)\�&��x   x   �!����%���JT�~���vν�H���8�`�j����И���Uþ@�ؾ���hG�����rG���@�ؾ�UþϘ�����]�j���8��H��vν�}���JT������x   x   `���_�	���'�S�X�����P���]���� �pH���q����nE���L�� ���u���n��������L��qE�������q�pH�� �b���O���������X��'�y�	�����x   x   ����'��_>�y6b�p+��4u���۽���O-%��RC�S2`�?�y�4����ꌾ%���ꌾ9���0�y�O2`��RC�G-%�����۽6u��r+���6b�Z_>���'����@��x   x   ~.T�joX��)b�ϓt�/c���q�������߽}�����"+�?T;��G�>M�,>M��G�>T;��"+���w���߽�����q��/c����t�*b��oX��.T��R���R�x   x   Vg��Ns��L���[������#�� 1��?s���@̽�?�����������՗�����������?��@̽Is�� 1���"�������[��G��Rs��&g���5�������5��x   x   ~Uν޾��]��da�����k��L������KC�� ��g���=丽�{���{��U丽m��� ��WC�����[���������Qa���]��޾��Uν�Pڽd��s�ཙPڽx   x   
2����T�ڽ����: �����y^��p�]�j��l��Vp��Wt���u��Wt�vVp��l�N�j��p�r^����% ������Y�ڽ���2��R�F �N#�&F ��R�x   x   l�8�� ����:�߽Z��Ip��F�o�91K���3���&�c ���"��c ���&���3�-1K�V�o�Ip��)Z��C�߽����� �y�8�2M�.	\�B�c�/�c�3	\�0M�x   x   ��j�DPH�Q%�ȥ�" ̽�,���j�X�3��%������ؼ�fѼs�ؼ���c%�j�3�Ңj��,�� ̽¥�G%�TPH���j�]ʄ�����֘�x����֘����dʄ�x   x   W���܎q�73C������{䥽�k���&�|���"��R4��y4��$#�������&��k��䥽����F3C�ڎq�R���g}������*�ľ o˾&o˾*�ľ����f}��x   x   ́��*�`�~+�����.m���,p��I ��ؼ*��ˌ�*����ؼ�I ��,p�m�������+��`�'ˁ����ƾO�߾+󾞝���������'+�M�߾��ƾx   x   =þ�/��%dy�96;��p��¸��*t�����FѼ�$���$��8GѼ����*t�
ø��p�66;� dy��/��%=þ��������������������#����x   x   k�ؾ�5�������F�l��Y����u�v��n�ؼ���Z�ؼp����u��Y���k���F����6��k�ؾ������_�'�o5�$Q>��_A�'Q>�o5�\�'�������x   x   j��<帾�׌��M�΀��Z��8,t��G �g�����G �7,t��Z��؀��M��׌�7帾`��a:�av%�2�;�U2N���[�̦b�Ʀb���[�\2N�3�;�^v%�^:�x   x   �-�Ar������
!M��m��Ÿ��.p��&�D���&��.p��Ÿ��m�!M�����Ar���-�x�d�1�(L�E�c�e v�����������_ v�@�c�(L�e�1��x�x   x   A���fs���ٌ���F��s�Fq����k��3��3���k�0q���s���F��ٌ�ms��>���ξ�A 9�}�W�uGt�C�������F���F������F��qGt�y�W�F 9�Ѿ�x   x   �0�踾����$<;�N���饽J�j��$K�C�j�饽M���!<;������踾�0󾵿��;��^���~������u��-۠�9i��*۠��u��������~��^��;����x   x   ���p;���my�	+��"�>1��=�o�B�o�21���"�+��my�t;�� ��4{�i"9��^�?��X���R��s��� ��! ��w����R��U��?���^�k"9�2{�x   x   \�ؾ�6���`����*̽.s���U�?s��*̽����`��6��\�ؾ�>���1�F�W���~�8��V���hӯ�H���3��H��iӯ�[���7����~�E�W���1��>�x   x   �FþA����?C�7��
c��*������c��8���?C�C����Fþ��:|%�.L�6Mt�?����T���ԯ�������������|ԯ��T��A���8Mt�.L�9|%���x   x   �����q��%��߽"'��*��-'���߽�%��q�����Ѹ�����;�P�c�B��Wy������mJ���	���Ŀ�	��lJ������Wy��B��O�c��;����и�x   x   ���VaH�M������O��]������S��WaH����i�ƾ��W�'�<N��*v�����!࠿�$��I7������G7���$��!࠿�����*v�<N�V�'���j�ƾx   x   ��j��� ��۽l��)���l���۽�� ���j�N����߾m ��y5�i�[�����L��To���%���L��Z���L���%��Oo���L�����k�[��y5�m ��߾G���x   x   P�8�Z���|n��Bc��Gc���n��R���Y�8��ׄ�K����>�)���]>�i�b�<���M��:⠿����ٯ�ٯ�����>⠿�M��;��f�b��]>�+���>�Q����ׄ�x   x   C�y���*����t�*��p���C��&M����)�ľ����k���mA��b��������W}��"Z������$Z��X}����������b��mA�k�����%�ľx���&M�x   x   qνz���)<b�/<b����qν�f�g$\�Q蘾'�˾������>`>���[�1v��������� ��� ���������1v���[�8`>�������/�˾Z蘾i$\��f�x   x   	|��>�X�Ok>�C�X��{���pڽ�\ �)d�?�����˾t���L���~5��BN�,�c�<Xt���~�lF����~�AXt�/�c��BN��~5�O��{�����˾1���'d��\ ��pڽx   x   �KT��'��'��KT�FM��&��q##��d��꘾_�ľ�E�V%��'���;��8L���W��^� ^���W��8L���;��'�X%��E�Z�ľ�꘾�d�y##�1��KM��x   x   ,����	�#����R�h�������^ �G)\����ܢ��q�߾l����� �%��1��/9�n�;��/9��1��%����f��r�߾墷����E)\��^ ����^�����R�x   x   �������9��?�R�pN��Wtڽk�{.M�|݄�������ƾ ��֤��H��������������H�Ѥ�"�澥�ƾ����|݄�{.M�k�xtڽpN��W�R�Z��x   x   2"׼�*��v��F��w������� ��")���V��ȃ����в��_ƾ�jվ��޾i⾺�޾�jվ�_ƾ�в�!���ȃ���V��")��� ����lw���F��v��*�x   x   # �z�.��P�I�<���o�����彨
���6��\�ݮ���g��0����������������"0���g��׮����\���6��
����f���@�����I�J����D �x   x   #i��z��1� 	R��b������Ƚ۟���)��s1�S�K��b���t�-����0����t�ͻb�P�K��s1��)�ʟ���Ƚ���b��.	R���1��z��h����x   x   V�E�]�I���Q��b��s|�$���mf��C�ʽt���	�9G���(�r3�R9�X9�r3���(�CG��	�g��K�ʽ�f������s|��b���Q���I�h�E���D�ѳD�x   x   �b�������U��f|�S���f��/��驢�Ph��Y˽�߽Z9�~���Lw��|���S9��߽�X˽Qh�������.���f��d��	f|��U�������b��>���^G��G���x   x   ~�����C���G_���s�dX|��U��L���Đ��|��v��7R��-R��%v���|���Đ�V���U���X|��s�O_��,��������󽽔ɽ�$Ͻ�$Ͻdɽx   x   �� ������ǽO�����bI|�+`��<O�O�G�=wF��|H�S�J�� L�7�J�~|H�HwF�A�G��<O�`�UI|����O���ǽ���� �����/�g���/����x   x   �)�����w��]�ʽؒ��?G��4/O��*��h�m��O����6�7򼃣������h��*�L/O�@G��쒢�c�ʽvw������)�G�;�g�I�)Q�Q�e�I�C�;�x   x   �V�s�6������YJ�����ݑG�^��ۼ���a����Č�뤔�������ۼ+^���G����OJ���������6��V�vFs�
ꄾv(��8���z(��ꄾ�Fs�x   x   Ե��+f\��V1��	�H5˽����;VF��������jm�59�F59�m�铭����UVF�����H5˽�	��V1�(f\�͵��n����H��lQ����������mQ���H��k���x   x   ������;�K�--���޽�_���UH��s�����]!9��7�M!9������s���UH��_����޽5-�4�K�������O+���!;p߾Y�� y�Q��u߾�!;L+��x   x   ǹ��PS����b�ƾ(���W��7�J�k�G���9��9�������6�J�&W����þ(���b�PS��ʹ��fvӾ�X��9�����:����X�dvӾx   x   Hƾ'��G�t��U3�ޞ���2���K�� ������l�ڄ��q ���K��2��Þ���U3�G�t�.��Hƾ��e	���I&�6\.��"1�6\.�I&����e	���x   x   mRվ�꨾����8�nL���3����J��o��3���w����o��
�J��3��uL���8����{꨾cRվ���<���+���<�N�H��6O�~6O�M�H���<�!�+�7�����x   x   ��޾�������A�8�����Y���VH����f�ۼt���VH�|Y��ˡ��D�8���������޾_	�/�"���:��P�`�`��Uk���n��Uk�Z�`��P���:�3�"�^	�x   x   ����$
���X3�Q�c���VF�WV�]V��VF��b��m��X3�&
���������q�)�ݐE�M_�Net��偿���������偿Tet�K_�ِE�r�)����x   x   ��޾����t�!�(�X�޽A���7�G��u*�(�G�I���T�޽�(���t�����޾���4,�`K�;�h��<��n������e7������n���<��?�h�^K�3,����x   x   �Wվ& ��-�b��3��=˽#��\*O�f*O����=˽�3�<�b�* ���Wվ�	�h�)��K���k�s鄿ـ��鞚�]j��aj��힚�׀��q鄿��k��K�g�)��	�x   x   hOƾ�Y����K�	� S��aI���`�mI���R��	���K��Y��kOƾd����"�H�E��h�:ꄿ�����(�������#�������(������:ꄿ�h�G�E���"�c��x   x   �²�i���b1�������LJ|�J|��������b1�m����²������:�w_��>�������)������?���?������)�������>��y_��:������x   x   ����u\�H�m�ʽ�%��Pp��%��k�ʽF��u\�����ӾHl	�$�+�$P�qlt�lq����������A��k尿A����������kq��qlt�$P�$�+�Hl	��Ӿx   x   �����6�����,[��c��%c��[��������6�����7���g�����<���`�[ꁿ2���An���&��%B��!B���&��Dn��2���[ꁿ��`���<����g��7��x   x   ��V��XȽ�����������eȽ	���V�/���71;�!��R&���H��`k������<��Io��Ϙ��$��՘��Ho���<�������`k���H��R&��!�=1;&���x   x   )�n�彠����s|��s|�����a��)��^s��W���(߾���g.��BO��
o�l�����������-���-���������n����
o��BO��g.���(߾�W���^s�x   x   `� �����Va���b�Va������e� � <�6����b��֝�}���/1�DO��ck��쁿�t��*���,���,����t���쁿�ck�DO��/1���ם��b��1����<�x   x   ���@���R�R�9��������L�I�b8���������}���i.���H�N�`�<tt��C���������C��7tt�Q�`���H��i.�|���������h8��M�I���x   x   �u���I�j�1��I��u��}2ɽsD��4Q�t���P�����k�QW&���<�,P�Z"_���h���k���h�^"_�,P���<�PW&�l���T���g����4Q�iD�o2ɽx   x   �F��������F��
��*DϽq��6Q�v:���f���.߾&�.����+���:���E�J(K�O(K���E���:���+�3��&��.߾�f��x:��6Q�x��4DϽ�
��x   x   �y��$��y���D��]��EϽ�F���I�����]���9;s�s	����|�"�R�)�C,�P�)�{�"�����s	�s��9;�]�������I��F�~EϽ�]����D�x   x   0�=0���O�D�����5ɽ ���<��is�篗�HB��L�ӾD��ݎ��	������	�ߎ�=��O�ӾLB��ᯗ��is��<���6ɽ���f�D�0��x   x   ��Ƽa�׼����3�8Cx��Ī�`u�/���?���k�Ւ��������v3����Ǿ�ʾ��Ǿv3��������ے����k���?�/�fu��Ī��Bx���3�~�V�׼x   x   ��׼�����987��o�������ͽ=J�1*#���D���e�"ˁ�C.����������������E.��+ˁ��e���D�;*#�;J���ͽ�����o�q87������׼x   x   ������"�k�>��g�e����Ѳ�ˣܽ�����5�?�I�f�Y���c�Gvg���c�o�Y�0�I�}5�#�������ܽ�Ѳ�l����g�y�>�:"�z��w����x   x   ��3��&7�S~>��_L�7c�+b����������P�ҽ��`[�+6�;���#��#�5��/6�c[���H�ҽ��������b��27c��_L�n~>��&7���3��2���2�x   x   rx��o��g��*c�N4e��o�1����w���H��{>��{@ý7ѽ`ڽk�ݽ`ڽ7ѽ�@ýx>���H���w������o�H4e��*c��g�Ւo�:x��w~��e���w~�x   x   ᩪ�𧝽l����T��c�o�MMb�:�]��a���k��y�f ��Z����󌽧�q���b ���y���k��a�S�]�MMb�x�o��T��t���⧝�詪����/��6��򞴽x   x   IP潵}ͽ����ɤ��n�����]���B���1��)�MP&���&�l(�Ŀ(�I(���&�QP&��)���1���B���]�]���Ҥ�������}ͽ]P�Vv�������tv��x   x   ,��4��ܽ@㳽@c��0�a���1�������Ѽ�x���j��&k���x����Ѽ�������1�3�a�Qc��C㳽�ܽ�4�*��(�}4�
;��	;�}4��(�x   x   `�?�#�g}���ҽ�-����k��)��������pz��I��:�q�I��pz�ԙ����)���k��-����ҽd}�##�f�?�؇Y�7�m���z��J��z�2�m��Y�x   x   �`k���D�4��^�q��r�y��2&��Ѽ�Tz�!A����������A�vUz�߈Ѽ�2&�b�y�s��"^�<����D�`k����+���9{��u&��t&��;{��)������x   x   ���we���4��C�|ý[惽��&�`M���fI�#����|������eI��M����&�W惽}ý�C���4�we��������η���Ǿ�?Ҿ��վ�?Ҿ��Ǿ�η����x   x   y쟾丁�N|I�"��ѽj���A�'�:��N�9����؛���9�^:��A�'�q����ѽ�M|I�渁�x쟾|��jؾ���Q���������S������jؾ
|��x   x   ���P��j�Y�{x��8ڽ-׌�Ҙ(�#9���XI�l"�qXI��8����(�5׌��8ڽxx�m�Y�T��	���aվ����R�	���
O�f��O���O�	�����hվx   x   ������c�6f#��iݽ�׌���'��H���8z�l9z��H����'��׌��iݽ<f#���c�����#X辬!��4�1*)��3��{9��{9��3�5*)��4��!�X�x   x   >�Ǿ퇛�OWg�Cg#�W;ڽp���'�&��Ѽ�����Ѽ�&�a���F;ڽHg#�DWg�퇛�I�Ǿ+��������'�@W:���H��CR��uU��CR���H�=W:���'����+���x   x   s�ʾማ���c�|{�~ѽ都L2&�V��W��`2&�都�ѽ�{���c�创�l�ʾ��55�k
1���G��>Z���g���n���n���g��>Z���G�h
1�35���x   x   ��Ǿ{��Y��!�#ýz�y�g)����_)�x�y�#ý�!� �Y�}򖾵�Ǿ���%T�c�5���O�3�f�+Ax��Ɓ�޷���Ɓ�&Ax�3�f���O�c�5�&T����x   x   T"�������I��I��%���k�w�1�}�1��k��%���I��I����L"�������6�m�5�$�R���l�#d��F@��G_��J_��H@��#d����l�$�R�o�5��6�����x   x   ����������4�;k�U5��K�a���B�T�a�L5��Dk���4���������_�K�t1�*�O��l��2���(���������􆓿�(���2���l�)�O�t1�O�_�x   x   ���I�e�G��ٝҽ�i����]���]��i��םҽD��R�e�����kվx&���'�/�G�(�f��e���)��(���?��B��*����)���e��)�f�0�G���'�v&�qվx   x   ������D�f��{ﳽZ����Ib�\���}ﳽe����D���������y���;��]:��DZ��Fx��B������-���[��-�������B���Fx��DZ��]:�;�z�������x   x   �rk��#�R�ܽI�����o���o�=���V�ܽ�#��rk�<&��Jwؾ��	�
2)���H���g�\ʁ��b��Ǻ�� ����ƺ���b��]ʁ���g���H�
2)���	�Cwؾ<&��x   x    �?��A��Ʋ�]���6e�]���Ʋ��A�'�?������ܷ����j'�m�3�~MR�V�n������c������秕������c������V�n�MR�p�3�g'���ܷ�{���x   x   J'���ͽ�����6c�w6c�������ͽI'���Y�ֵ���Ⱦ����7Y���9��U�лn��ˁ�;E��6-��4-��9E���ˁ�ӻn��U���9�7Y������Ⱦص����Y�x   x   �k潿���$�g�DgL�0�g�ǹ���k�W'(���m�ꊡ�nRҾ�����ć9�&PR�	�g�Mx��i���7���i��Mx��g�$PR�Ň9������sRҾ芡���m�P'(�x   x   ���p�o���>�Ȍ>�K�o�������R�4���z��7����վ��@[���3��I��KZ���f�9m�<m���f��KZ��I���3�A[�����վ�7����z�S�4�����x   x   �?x�~:7��"��:7��?x�ʸ��Z���";�ri�9��UUҾ����T+�z7)��d:��G�n�O���R�j�O��G��d:�x7)�P+�����_UҾ9��`i��";�T������x   x   ��3�������3���~�Q���(��#;�D�z�j���Ⱦ����	�B��'�m1�� 6�� 6�o1��'��A� �	����vȾe���@�z��#;��(�Y��ܝ~�x   x   $��(�M���2��y��~��F��P�4���m�K���N䷾��ؾ����y.����A��_��A���{.�������ؾT䷾O�����m�W�4�5�����y��}�2�x   x   �׼�׼'��9�2���~�廴�����-(�T�Y�v����/������,վ"p���� ��������%p��,վ�����/��s���V�Y��-(�
��� ���~�L�2�T��x   x   ȷ�������6�w��Z�+����]ɽ���^Z'��^M���s�ʋ�%W���U���殾B|���殾�U�� W��ʋ���s��^M�YZ'����^ɽ<�����Z�"w�h6Ｆ���x   x   n�����ռ�C �)Z"��AS��]��0������+��7+���G�mCb�S	x�˃��ׇ��ׇ�˃�P	x�}Cb���G��7+�,���5����]��BS�BZ"��C ���ռ<���x   x   �!�`= ���(��1L���{��2��B!��X5��	�P<��"/��-=��"F�c6I��"F��-=��"/�K<��	�g5�?!���2����{��1L���(��
�S= ��!�M��x   x   ac��J"�*�(���4��
H�G�d�3���c��v���U�ѽ���q� �	�HP�GP�	�p� ����i�ѽs���vc��3��G�d�H�~�4�F�(�K"�Mc�)a�a�x   x   �Z�'S��L�= H��1I��fQ�vHa�D>x�y'���;������c��g(���ݽ�k(���c��*����;��i'��O>x�zHa�gQ��1I�E H�L��&S��Z���_���a���_�x   x   ����rI����{�hid�B[Q���D�.�?���A�:YI�k,T���_���h��n��n���h���_�X,T�;YI���A�>�?���D�V[Q�sid���{�bI�������:���㢽�㢽�:��x   x   �=ɽ����$��!���0a���?���&���������	�Gb	��	�l@
��	�Qb	���	���������&���?��0a�!���������=ɽ��ڽ�,潗!꽟,���ڽx   x   ����������J���x�/�A�7���������A楼�𕼫ӎ��ӎ���\楼������G��@�A��x��J�����������_��{o�##�##�to�a��x   x   �@'�f����ix��$��(9I�a�����p����13��������^13�C���>���o��69I���hx����h���@'��=��O���Z���^���Z��O�	�=�x   x   �@M�+�]����ѽ����T���	��ȥ��3��q���������r��<3��ȥ���	�]T����ζѽ]��+��@M���l�ř��H��A��<��K��ƙ����l�x   x   �~s���G��"�Ģ뽙s��Y_�mC	��ʕ��W�)���G���W��ʕ�^C	�Y_��s������"���G� s�E����Ǡ�����1�����/�������Ǡ�G���x   x   跋�J#b��/�{� �
B����h���	������b��b��c��c������	���h�B��t� ��/�R#b�ⷋ�Υ�~���.5ѾnB߾j��r��oB߾*5Ѿ~���Υ�x   x   D����w��=�c�������m�
�[���qK�^9���J�E����
���m����c���=���w� D��.����"ؾ������	��7��	��������"ؾ0���x   x   �B��9����F��9�������m���	��ŕ���2�%�2�ƕ���	���m������9��F�5����B��\�˾���JM��_�|����"���"�}���_�LM����U�˾x   x   �Ӯ�8Ǉ�I��:�����h��C	�￥�ፂ�����zC	���h����:�I�9Ǉ��Ӯ���׾b$ ��
��b#�	0��8���:��8�0��b#��
�e$ �þ׾x   x   "j��ȇ�/	F� ��,F��s]_���	����������	��]_�7F����.	F�ȇ�j��J�ݾz���U���.��>���J�N�P�K�P���J��>���.��U�v��L�ݾx   x   �ծ������=��� �By��H	T����������1	T�:y���� ��=������ծ���ݾ�{�����6�\�I���X��Nb�F�e��Nb���X�Z�I��6�����{���ݾx   x   �F����w�c/����%��2=I�*��*��?=I��%����j/���w��F����׾�����ܗ8�5O��a���n�)�u�+�u���n�!�a�5O�ؗ8��������׾x   x   �I���-b�
+��ѽF��m�A� �&�j�A�?���ѽ+�z-b��I����˾_' ��X�� 6�_O�8�d�p�u��*�����*��o�u�6�d�`O�� 6��X�b' �|�˾x   x   ����U�G�������i%x��?��?�n%x�������Z�G�����-���3������.�I���a�֜u��򁿦���������֜u���a���I���.���1��2���x   x   ��s�A)+� �+U���8a��D��8a�/U�� �C)+���s�Pץ�`-ؾ�R�7h#�~?���X��o�,��m��� ���m���,���o���X�?�9h#��R�a-ؾOץ�x   x   �PM�\	�����)��X`Q�\`Q��)�����\	��PM�D���*������f�0�܇J�$Ub���u�[��8���8���[����u�$Ub�އJ�0��f����%���D���x   x   AP'�����(��Cwd��3I�Pwd��(�����EP'�
�l��Ӡ�=CѾA�����f8���P�.�e�L�u��-���􁿊-��K�u�,�e���P�d8����@��@CѾ�Ӡ���l�x   x   ���������{�F
H�2
H���{����������=�ȥ��J���R߾�	�%�"���:��P��Wb�#o���u���u�"o��Wb��P���:�&�"��	��R߾D��ɥ���=�x   x   �Uɽ�X��S/L��4�^/L��X���Uɽ>���O�'��r������A�.�"��8���J�ɾX�l�a�Y�d�j�a�˾X���J��8�-�"��A�æ�y��'���O�6��x   x   �����>S���(���(��>S���ڽ݂���Z�� ���1��O��r	����j0�W
?��I�!O�!O��I�U
?�k0����t	�N�澷1��� ����Z�߂�,�ڽx   x   �Z�\"�"�)\"��Z�4Q��\L�c8#���^��!����HW߾���Mk�Wn#�'�.��)6�١8��)6�'�.�Xn#�Lk����DW߾	���!����^�d8#�TL�%Q��x   x   �w��H ��H ��w��`�2����C꽕9#���Z�(*��2��YJѾE���X�_�4a�f��f��4a�`��X�I��`JѾ.��$*����Z��9#��C�=����`�x   x   ;���ռ�;�Nw�`!b�9����O�U��>�O������ڠ�T����8ؾM�/ �Y����[���/ �L���8ؾO����ڠ�����G�O�_���O�;���+!b�?w�x   x   ӑ����������v�Q `��S��^�ڽ�����=�9�l������᥾�����˾��׾�޾޾��׾��˾����᥾����>�l���=����O�ڽ�S��m `�w���x   x   ����/���м�	�>�;�������H^�E�=�.��WO�a8n�m���gᎾ	n�����n��kᎾk���V8n�	XO�<�.�E�C^�$������4�;��	��м�/��x   x   �(��������޼�^���5� �l��B����½Dd�e���)�7Y@��S�b`��Yg��Yg�b`��S�AY@���)��e�2d񽹼½�B����l���5��^�-�޼ᕺ�r(��x   x   �м�޼����D����/���W��@��?]��@ŽZD�>?��p�Ec ��(�h�*��(�Oc ��p�3?�ED�cŽE]���@����W�Ѻ/�R��������޼_мnI˼x   x   b�	��Q��������,�w�C��c��̄�����kc��Gǽ��ٽ�T�݂�ւ��T罰�ٽ;ǽ�c�������̄��c���C��,��������Q�T�	�U��*��x   x   \�;�ѡ5��/��,�Ѭ,�� 3�l�?��0R�Ei�(䀽ȱ��s�����V��%���s��ڱ��$䀽"i��0R���?�� 3���,��,�+�/���5�r�;�o@�B�o@�x   x   ~��j�l��W�+�C���2�B�'�Je"��#���(���0���9���@��E��E�r�@���9���0���(��#�Te"� �'���2�L�C��W�Z�l�����C���3���3���C��x   x   ތ���*���,��3�b�E�?�z["�\e����|��4p�;�޼��޼��޼�޼r�޼�o�ȱ���e��["�h�?�7�b��,��~*������ef���ĽCiǽ�Ľ|f��x   x   �:�A�½�B�����mR��#�M	���¼$S��$����Ve���W���W�GVe�0���+S����¼f	���#�hR������B��a�½�:�Rq��0����
���
�,��Xq��x   x   Y/��=�u�Ľc�����h�`o(����D����F�����^���ߍ�W^��z�����F��D����jo(���h�l�����Ľ�=�Q/��`!�!�0��6:���=��6:��0��`!�x   x   ��.��N���OD��h̀�ޤ0��C�Ќ��Q���H�%��^���5��t�%����������CἭ�0�ò�gD�����N���.��I�u)`�cpp�m�x�\�x�ipp�})`��I�x   x   ";O�?�)��)�[�ƽ�����x9�x�޼�e�s��	8���4�:�2������e�~�޼�x9����P�ƽ�)�C�)�/;O�a�r�R)���b���'���џ��'���b��V)��j�r�x   x   n��=@�MY�>�ٽPV����@�[�޼szW�������燍��zW�|�޼��@�EV��1�ٽQY��=@�n�������������.Wž4Wž�����������x   x   s���R�K �@.罐���D���޼�wW�� ��d%�v����wW���޼��D���F.�&K ��R� s��S���d���ZϾ$����ר��$�\Ͼa���P���x   x   �Ў�
E`�e�'�Y\�4����D���޼�e��v���w��e���޼��D�0��P\�]�'�E`��Ў��M����̾;�{����B��k��k��B�r���>辶�̾�M��x   x   �]���=g��*��]�yĜ��@�V�޼������F�b���%�޼�@�xĜ��]��*��=g��]��]ĸ�(�۾�[�� 2�?�z���+ �y��?�2�}[��,�۾dĸ�x   x   j���?g���'��2��Y��T|9��A�x7���7���A�i|9��Y���2罉�'��>g�e����0��4J��V�����#�Y�-�D�2�A�2�Z�-���#����V�,J��0��x   x   y_��SI`�KO ��ٽ������0����¼���h�0������ٽLO �RI`�_��2�����	��C�g�,�@�9���A�-ZD���A�=�9�c�,��C�	����2��x   x   TԎ���R�_��ǽ�р�Nr(���������lr(��р��ǽ_���R�RԎ��Ǹ��L��	��`�s1��A�^9L�|R�{R�\9L��A�	s1��`��	��L徽Ǹ�x   x   x��]F@�l0��M����h�##��]�#���h��M��p0�^F@�x��/S��Y�۾Y�rE�t1��C�\�Q�W�Z���]�X�Z�Z�Q�߫C�t1�vE�Y�V�۾-S��x   x   2%n�2�)�l,�ϋ��=R��Z"��Z"�6R�ۋ��o,�/�)�/%n�?���	�̾�b��N�I�,��A���Q��]���c���c� �]���Q��A�G�,�K��b���̾@���x   x   �HO�EY� �Ľ�����?���'� �?������ĽFY��HO����g�����6���#�a�9��<L�ʩZ���c�}�f���c�ǩZ��<L�`�9���#��6���i�����x   x   \�.��Q�8P���c���2���2��c�0P���Q�\�.��
s�/���ϾW���C�1�-��A�2
R�}�]�D�c�E�c��]�2
R��A�4�-�C�Q����Ͼ.���
s�x   x   {<�د½}8��ĬC��,�άC�8���½u<�6�I��3������v1��I����P�2��`D�kR�S�Z��]�O�Z�lR��`D�N�2�����I�|1������3��2�I�x   x   �Rང:���W�,�
,��W�x:���R��p!�>`�.o�����.�t��3 �`�2�f�A�Z@L�`�Q�e�Q�\@L�c�A�`�2��3 �t�(����-o��>`��p!�x   x   ���>�l���/������/�c�l���������0��p��5��gž���t����S�-�Đ9��A���C��A�Ő9�U�-�����t���gž�5���p� �0����x   x   �	���5�s��{����5��	��E~�����1L:��y�៾^hž6뾈L��
���#�s�,�X{1�X{1�t�,���#��
��L�9�^hž៾�y�'L:����M~��x   x   ��;�G`�����c`���;�MV���)Ľ��
�ؤ=�iy��7�����c7�m���<����L�5i� M���<�p���`7�����7��ty��=���
��)ĽBV��x   x   ��	���޼^�޼��	���@�?H���ǽ��
��N:�Z�p�cs�� ���"ϾP"辒o���`�O	�L	��`��o��M"��"Ͼ ��gs��V�p��N:���
��ǽOH��׊@�x   x   �м�Xм��f<B�"I���,Ľ���R�0�QF`��9����k��;�̾��۾�\復��]徕�۾5�̾p�����9��IF`�a�0�����,Ľ&I��4<B���x   x   /3��3��_˼���&�@��X������0���x!���I��s����Q���4`���ָ�rB��nB���ָ�7`��T�������s���I�x!���������X��4�@����Q_˼x   x   6ǅ�FX�� ������U����U��ώ��,����뽇����+�C�E��B\�l�m���x���|���x�t�m��B\�;�E���+������뽫,���ώ���U�l����輾���=X��x   x   jR���ݞ������7��d	F��"�����I�ǽ���ޠ��P���.�=:�B�?�R�?�@:���.��P���~��-�ǽ�����"�R	F�6��P��� ޞ�UR��x   x   /������oӼ���դ���4�u�]������������(ܽ-@��Ą���
�����
�ʄ�F@���'ܽ�����������d�]���4�ڤ����"oӼr�����'���x   x   G��&��V���<��w��#�F=��,\����#O���	���@���d��CHĽ7HĽ�d��q@���	��EO������,\�<=�$�#��w��<�h����B���>缠>�x   x   (��}����yp����j�;�N�-�I	@���S���f�dv�x^��-���^��	dv���f���S�7	@�J�-�6;��j����p� ��_��H��}�!���"���!�x   x   �U���E��k4�:�#��b�7i��l��D���	�P����S�ˀ����S���^���	�E��l��h��b�F�#��k4���E�%�U���a�\h�\h���a�x   x   w���H�~���]�7�<�p*��d����_�̼�����G���尼���0������5氼CG��7���x�̼)���d��*�;�<�z�]�7�~�{���h������ƥ�p��u��x   x   ����~���s��\
\�\�-�85�ó̼RZ��'�s�}0F�,+�ó�����+�k0F��s�Z��ҳ̼P5�K�-�-
\��s���~�����,�ν5޽?>�R>�5޽(�νx   x   {��J�ǽi���Jc���?�>�	�싼�.�s�ϔ������>�R��>����M��N�s����D�	�{�?�fc�����6�ǽn�뽻���b�Cv�b>�Gv��b����x   x   >��ы�ۿ�g5��d�S�3���"�� F��v���,9�Ĺ:ƹ:_/9��v���F��"����n�S�x5���ڿ�̋�D���''��:�K�G�2�N�"�N�M�G��:��''�x   x   ��+����*ܽ�죽#�f�������*�!j>��%�:�s9;�%�:j>���*�������=�f��죽)ܽ�����+�ƿI�qd���x�Ղ����Ղ���x�ud�пI�x   x   ��E��9�f��Z!��G4v��0�zۯ�u�W���`�:�^�:��&u��ۯ��0�,4v�T!��f���9��E��ek�6솾D4��l����������l��C4��2솾�ek�x   x   \'\���.��p��D���E��]��ǯ�tr�D>�a�7��B>��r��ǯ�]�F���D���p���.�V'\�愾Ea��.��au���ľ��Ǿ�ľgu��1��Da���儾x   x   Q�m���9���
�/(Ľ����]��ۯ���*�2M���M����*��ۯ��]����(Ľ��
���9�]�m�8d��R���;¾<վͽ⾖�龟��ѽ�<վ�;¾X��7d��x   x   6�x�a�?�C��c)Ľ�G���2�����D�E�ct���E�_����2��G��\)ĽV��e�?�3�x��D���췾K{Ӿ�*�zc���o��e��o�{c���*�D{Ӿ�췾�D��x   x   z|���?�~�
�PH���9v�X�� ����s�؞s�` ��e���9v�ZH��y�
���?�z|�����] ��ե߾����\y	�x��U��U��y��\y	�����ץ߾W ������x   x   M�x�u:�t��&����f���G���I��"��������f��&��t�t:�W�x��ើ(�¾���y/�E����h"�{�$�!h"����A�z/����,�¾�ើx   x   b�m�K�.�#���󣽖�S�K�	�8�̼-�̼o�	���S����"��O�.�f�m��G������徉����+"��=+�g0�c0��=+�2"��������徨���G��x   x   �/\��@�Zܽ9=����?�16����(6���?�'=��qܽ�@��/\��h��񷾺�߾�0�R���($�^�/�2&7�!�9�8&7�\�/��($�T���0���߾�𷾼h��x   x   ,�E���翽�r�S�-��c��c�F�-��r�翽ޓ�*�E��넾�����Ӿ�������"�U�/���9���>���>���9�Y�/��"���������Ӿ����넾x   x   ��+����t��4\��/��e��/�6\�n�������+�Bsk��h���C¾�2�;}	���\@+�6(7�Φ>�6A�ͦ>�5(7�\@+���<}	��2��C¾�h��=sk�x   x   �����ǽ�~���<��e��e��<��~����ǽ���,�I��􆾮��"Fվ�m��`���l"�L0�7�9�ݧ>��>�:�9�I0��l"�d���m��Fվ�����7�I�x   x   =��ݍ��t�]���#�����#�z�]��&���5'�d��>����������u�=����$�K0�P*7��9�I*7�L0��$�;���u����À���>��d��5'�x   x   #����r{4�:w�Aw�b{4�n�
#��!��:�x�x�x���ľP���l�!���n"�NC+�V�/�[�/�RC+��n"� ���l�U����ľx���x�:���x   x   ʎ�;F����@���^F�ʎ��Ͻ�r��G����� ͤ��Ǿ���}w��������"��.$��"������zw�����Ǿͤ�����"�G��r��Ͻx   x   ��U�������������U���;P޽��*�N����#Τ���ľ ���s��c�	���u��t����d�	��s�� �⾑�ľ%Τ����!�N����DP޽��x   x   |�����zӼ&�����a����6\潟Q���N��₾O{�������Lվ�;�r���M7����Q7�l����;��Lվ����K{���₾��N��Q�;\潤����a�x   x   �����������[�!��}h��ޥ��]�V����G���x��C������L¾G�Ӿ]�߾[ �S �Y�߾U�Ӿ�L¾����C����x���G�C���]潬ޥ�~h�h�!�x   x   ���Y瞼I����]���"�]h����&U޽�v��$:�'d�^���_q���'�����F��$�¾N������'��dq��c����&d��$:�
w�2U޽���gh���"��]�x   x   ;[��0[��ʬ�o]缉�!���a�k��mϽ)���>'��I���k�1����s��@T����AT���s��4���z�k��I��>'�#��gϽ`����a���!��]�Iʬ�x   x   0�_���p����K������.��h�������:��%�
�d��I&2��v@��I�ƨL��I��v@�P&2�a���
�5��ك������|h���.�6���K������p�x   x   �p��?��CҜ�o�üϬ��8�!��ZO�fӂ��s��{½f�⽫t ���y1�{�����~1����t �}�⽇½�s��Zӂ��ZO�G�!�ɬ��:�üKҜ��?���p�x   x   �����ʜ���H�ʼ�X�d��L4��Z[�w���R���s*���NŽ�:ս�o߽[���o߽�:ս�NŽm*��9��������Z[��L4��d��X�T�ʼ���ʜ�����_���x   x   )5���üp�ʼf�׼���w��o���1���M�Ak�ݲ���ˏ�����u\��i\�������ˏ�ڲ��&Ak���M���1��o��w��켁�׼r�ʼ�ü.5��_���G���x   x   <{������B�#��gl켇)�n� �R/�mE��)�h8�=�D���L���O���L�P�D�h8�	�)�vE�M/�� ��)�l�5��_B����S{����'�����x   x   `�.�R�!�fR�k�m�����ؼFq׼]*ܼL��9�����i���Y�������;���=*ܼLq׼��ؼ��f��j�_R�y�!�^�.��S8���=���=�T8�x   x   ��g��:O�924��[�� ���ؼH$��2����O���V������+S���
��_S�������V���O��9���I$����ؼ� ��[�T24��:O�t�g�L�{��d��]����d��S�{�x   x   ��������7[�4�1�?��W׼`����9t�޷9��a�c���g߻g߻b���a�ѷ9��9t�]����W׼/�'�1��7[��������(��� ﳽ�p���p��ﳽ���x   x   �f��Z���}����M�+� ܼ:��X�9�$һ�L��6���[%��9���L��һY�9��9��ܼ$+��M��}���Y���f��LؽF������c������T��Lؽx   x   �z���������k�k�)�ՙ伺8��;?���K��k:�;�;l:��K��>��8��˙�k�)��k���������z齄��u���!�$d'�d'���!��u���x   x   ��
����u������BD8��a�뀈�����n����;��h;��;p��m�����b�ED8�~��������⽌�
��#��8�gwI�G2T�^�W�O2T�awI��8� #�x   x   ����a �o/Ž������D������+��� ߻4k#���;��;�h#� ߻�+��S�����D�����i/Ž�a ����>���Z�[r�q���� ��� ��r���#[r���Z��>�x   x   �2��ս되�$�L�ql��↼��޻�/���:~-���޻z↼dl��Q�L��	ս ��2�ۂW��z��׌��ɘ�\��n���\���ɘ��׌��z�҂W�x   x   �_@����N߽yB��jtO�jm���+������O�K��K�]����+��mm��ctO�iB���N߽���_@��l�]E���o���1���e��&8��-8��f���1���o��`E���l�x   x   PuI����h��lC����L����F���H2�t�ѻ2�+���.�����L�hC��������FuI�>�z�h땾[Ȭ�s���Ͼeپ�Yܾ[پ�Ͼs��VȬ�f땾D�z�x   x   ��L����Q߽̓���D��e�D6��7�9�D�9�u6��f��D�ѓ���Q߽����L��2��y����궾�bξÄ���J��M���﾿���bξ�궾u����2��x   x   �wI�� ��ս����I8�(�伎5���t��5��ܝ�J8�����ս� ��wI��3���r)���׾�!����g��J��g������!��׾u)����3��x   x   |d@��	�(7Ž���ʉ)��ܼ����֓��	ܼډ)����7Ž�	��d@���z�a����*���ھ����H�!����������M������ھ�*��^�����z�x   x   �2��g �y���#k�q1��X׼���X׼m1��#k�����g ��2�l���f ׾������*u��x�c���x�)u��������l ׾��l�x   x   D��W��(���
�M�� ���ؼ��ؼ� �"�M�+���C��B��z�W��J���ͬ��gξ�%����u�rv�I��F��pv��u����%gξ�ͬ��J��v�W�x   x   ��
��½6���<�1�� �,�� �:�1�4����½��
��>���z��v���y��5��y���u��;z�&��U��&��;z�u��v���6���y���v����z���>�x   x   !��Ig��_I[�"e�!�� �7e�JI[�Kg��0�齶+#���Z��ߌ�:��y�Ͼ �sk�ܣ���������٣�rk��z�Ͼ:���ߌ���Z��+#�x   x   =x���ʂ�lA4�Hr��m�Jr�iA4��ʂ�,x���z�8�	lr�+Ә��o��{#پ��\O�����{� y��{����`O���s#پ�o��/Ә�	lr�t�8��x   x   �����OO��^������켹^��OO������aؽ���o�I�J����f���C��weܾ���m���>y�Cy���m����|eܾ�C���f��I���v�I�~���aؽx   x   	h��!��U��׼�U򼘴!��h�������ԡ!��ET����� ���D��$&پXﾅ�����U��������[�&&پ�D��~ ������ET�١!�������x   x   ã.�+���t�ʼj�ʼ�����.���{��������v'���W����i���s����Ͼ��$.�������%.��ᾮ�Ͼ�s��i�������W�v'����������{�x   x   ���W�üt���{�ü����l8��v������3���<w'��HT����Iט��?��8����pξ�*׾�#ھ�*׾�pξ2����?��Nט������HT�=w'�M��������v���l8�x   x   �L��؜��ל�tL�� ����=�w������X���g�!�?�I��tr�\匾�}��z֬����i6��c6��|����֬��}��W匾�tr�K�I�n�!�B������k�����=�"��x   x   zŒ�<G���Œ��������=��x�������� ����8��Z���z�S�������������������S����z���Z���8����������x���=�������x   x   w�p�q�p�����<����p8��|�C���skؽ?#�m5#�}�>�ϛW�G1l���z�?��
?����z�B1l�ԛW�{�>�p5#�@#�fkؽI����|�p8�
��I�����x   x   �7���D�g�n�V|��4м��/^8�kln�N)��uɷ�Aڽ�@���%�W��k��:!�f��Y���%�A���@ڽlɷ�`)��vln�)^8���+4м_|����n���D�x   x   E�D��W��~�'���Wɼ$���$��N�0O~�d���������ɽ�xݽf���S��S�k���xݽ��ɽ����v���2O~���N���$�$��Wɼ#���~��W�@�D�x   x   �n���~����ӓ���h¼b$����*-�0O�ۮr��Պ�ℚ� ��쮽F����쮽��鄚��Պ�ʮr�O��*-��t$�ah¼ϓ�����x�~�B�n�;�i�x   x   �j��l��	���O����t��[lԼ���4��!��28�C�M���`��Pn���u���u��Pn���`�@�M��28��!��4����lԼt������
���j���j���x���x��x   x   �м�?ɼW¼(k���c��W���sh˼�ܼ�-�98��n������#!����!���n�+8��-�ܼ`h˼c���&d��(k���V¼�?ɼ�м�
ռb�ּ�
ռx   x   �k����>XԼ����I�����ߧ�ܚ���w���f���_��3���G����_���f��x��嚪��ާ�����I������WԼ�� �wk��6��e��e��6�x   x   �A8���$���+��mS˼����􏼹Rz���a��S���K��H���G�T�H�	�K��S�\�a��Rz�������PS˼6��<����$��A8�H�`PR���U�vPR��H�x   x   �Gn���N�a-�����ۼ˧�@z�8�R���&ͻ�Ԥ�R푻LԤ��&ͻa��p8��?z��ʧ���ۼ�]-�l�N��Gn�����S���y���y��S�����x   x   ����&~�	�N�u�!�q�)~���va�Ƈ�+���VǺe'(8�:J�'8�Ǻ9�������va�;~����z�!���N��&~����Ɣ��<Ⱥ�[,Žl�ȽQ,ŽNȺ�ɔ��x   x   `����p����r�;8�L��S����R�h�̻��ƺ�;�:bqC;nrC;�=�:ݿƺo�̻��R��S��B�8�~�r��p��^���ŶԽ*&�7���	�	�5���&�ֶԽx   x   "ڽ�ݱ������M��R�s=����K�T���
O<8L�C;,Q�;?�C;�<8(���ЉK�}=���R���M�1����ݱ�"ڽ�l �P�������'�x~*���'����O���l �x   x   	��}ɽ/l��p`����3��zkH�M���6�:-�C;�C;]�:ؚ���kH�3�����p`�)l��}ɽ
��H"�$�,�>�?��M�'T��&T��M�E�?��,�F"�x   x   ���Yݽ6ئ��'n����=����G�������B8W��: �B8���3�G�=�������'n�3ئ��Yݽ���)�EQF��_��\r���~��e����~��\r��_�NQF���)�x   x   �o�ذ��Ү��lu�� �����jH����{KƺiLƺ����jH������ ��lu��Ү����o��d:��\��{{�'���B���R��R��E���(����{{�
�\��d:�x   x   >���4�
���?nu�b���4���K���̻�͊���̻ՇK�5��w��Anu�����4�6��'F�"�m�#^��lX��s����i������i��u���lX��"^���m�~'F�x   x   �(!��6�ծ�,,n���2@����R�w��v���R�T@����),n�ծ��6�(!�]JL���x�8���U����O��	Y��Xž\ž
Y��}O��X���;�����x�YJL�x   x   G�����ܦ��v`�W��V���na���7��na��V��W��v`��ܦ����E���KL�7G|�jޕ��֫�����;:
־)پ<
־�; ����֫�iޕ�>G|��KL�x   x   �s� aݽ,r��$�M� $�)���*3z�*3z�1���#$�,�M�r���`ݽ�s�I+F���x�Qߕ�xE��$�þ?�վ���^�^����B�վ(�þ{E��Pߕ���x�H+F�x   x   ��0�ɽ3Ɗ��8��7˧��돼˧�:�8�8Ɗ�<�ɽ��j:��m�ܜ���ث�D�þ�xؾs� ��;��)��r辞xؾC�þ�ث�ޜ���m��j:�x   x   -,��/豽f�r�ʏ!��ۼX���������ۼˏ!�q�r�'豽*,��w�)�a�\�Ub��<���N�����վ���$��'���#����$���辬�վN���<���Sb��`�\�w�)�x   x   L0ڽP{����N��'�&Y˼ E��Y˼�'���N�N{��P0ڽ+�`[F���{��]���T���;���������jC����������ᾄ;�T���]����{�c[F�+�x   x   �����;~��-�]��>����������-�~;~������u �K�,��#_�񇊾[����_��S־Hc��?�����������?��Cc�T־�_��X��������#_�G�,��u �x   x   / ��4�N����cԼ�d��cԼ���@�N�/ ����Խ���Ǘ?�*lr�[����q��[ž�%پ�d辠��")�����d辟%پ[ž�q��Y���#lr�Ǘ?������Խx   x   `n��$���2s��Ds������$�`n����� <��j"M�*�~�O[��J���ž�־���"� "辮���־�žG��P[��.�~�o"M��<����x   x   �V8�v��e¼݋���e¼~��V8�ݝ��(ܺ������'��8T��o��P\���s��>c��y;�վ?�ؾ�վu;>c���s��P\���o���8T���'�����8ܺ�ܝ��x   x   <|��Tɼ���������Tɼ5|��)H��d���BŽ5�X�*�;:T���~�I�������bZ��M�����þ��þN���gZ������E�����~�=:T�_�*�8��BŽ�d���)H�x   x   �1м�����������1мHJ�1lR�������Ƚ6�p�'��&M��rr������c������t᫾4O��y᫾�����c�������rr��&M�i�'�3���Ƚ����PlR�CJ�x   x   }��J�~�F�~�}���'ռ,{�{�U������EŽS����	���?��,_���{��i��g����蕾�蕾f����i����{��,_���?��	�]����EŽ����c�U�{��'ռx   x   ��n�طW���n�ь��(�ּ�{�3oR��g���ẽ�D�1���,��fF��\�5�m��x�_[|��x�>�m��\��fF��,�4���D��ẽ�g��<oR� |�M�ּˌ��x   x   ��D���D�u�i�����#)ռ�L�#/H�����h���R�Խ�} �5��*�Ly:��;F�^L�^L��;F�Ay:��*�5��} �J�Խ`���â��/H��L�	)ռ�����i�x   x   +d����>�7�v������9ڼ%K�KE8�Og������%���G��|ֽt���������u��|ֽ�G���%������Sg�XE8�)K�o9ڼ~���0�v�:�>���x   x   �	�Ш,���J��Nz��]��h�ɼϫ��6���vC��i�9��r��'#������ҹ��ҹ����0#��g��0��(�i��vC�&������t�ɼ�]���Nz���J���,��	�x   x   �>���J���`��"������P��y�ݼ	l������9���S�\�k�kr~�=E��9[��IE��^r~�V�k���S���9�e���k���ݼ�P������"��{�`���J���>��:�x   x   �zv�o9z����$f�����H���\x���Q׼�2���o����,�*�I�4�#u:�$u:�G�4�0�*�����o��2���Q׼Xx��������Bf�����l9z��zv��u��u�x   x   �ޣ�BK���������l���┼����觼�=���Jȼ��ؼ��{�����_���漆�ؼ�Jȼ�=���觼����┼m��y��k��cK���ޣ�/է��C��:է�x   x   �ڼ��ɼ�:���夼�ڔ�����8b��A�}�x������Y��`p���̎��̎�hp��qY�� �������}�&b��'����ڔ��夼�:����ɼ�ڼ�`������켾`�x   x   �5�z����rݼ`�����GZ����X��9�U�$�6��\������!��U�C��#�$���9� �X�IZ��d��`���rݼt����5�H���#�UO&�7�#�<��x   x   C)8�H���V�*0׼;Ч�Xa}�j�9��}�=X�����yE��P%��O%��E�(��RX��~�\�9��`}�8Ч�V0׼�V�3��J)8�xM��-\��)d��)d��-\�zM�x   x   ��f��WC�e������� ��V�$��?��x� ������*�:L8�:(�:󠃹ɛ ��?��;�$�6��F�����G���WC���f��Y��叽�<����$叽�Y��x   x   C錽��i�9��V�T$ȼR���'���탻Wu��,�;L3\;�3\;�;-t��=6��[���=$ȼ�V�؁9���i�9錽U���:����ý�˽�˽��ý�:��U��x   x   ��~����S�����ؼ�9�����ĭD�˩�:hM\;ZL�;SM\;槅:k�D�����9���ؼ�����S�t�������Ľ�l߽-D��b� ���Y� �5D���l߽��Ľx   x   u-����~k�ӓ*�@]��M��1����$�z׻:�]\;@]\;Qػ:�$�E���M��?]�ؓ*��~k��}-��J*潕��?�����U#��U#����?����L*�x   x   W`ֽI���J~���4�3x�.�����@�$��ԅ:��;Յ:��$����3���.x���4��J~�L��^`ֽ|R��b�m�+�F�:��sD�t�G��sD�@�:�j�+��b�~R�x   x   ��v���R1���U:����Ʃ��w���D�K ������@�D�|��������U:�Y1��{������.�)���A��V��`d�l�k�e�k��`d�V��A�)�)��x   x   ���ʺ���G���V:��z�7O������ۃ�;R �B܃����>O���z��V:��G����������!��7��.T��rm�u}�������Ĉ�����u}���rm��.T��7��!�x   x   ��������3��&�4�8b�k;��J���$��Q$��J��;��$b�"�4�3�������������΋?�f)a��v�3(�����≙�≙����3(���v�g)a�ҋ?����x   x   �������fQ~��*���ؼ>���V�$��j�m�$�;�����ؼ�*�hQ~� �������IuB�A�g��f���e��I韾2&��2���1&��K韾�e���f��=�g�GuB����x   x    �������k���x+ȼ�����9�Ð9����k+ȼ����k�������$�8�?���g�9V��m����Ŧ�ະ��ൾ�ൾẰ��Ŧ�m���>V����g�2�?��$�x   x   �hֽ����c�S��]�%���`}��{X��`}�6%���]�W�S������hֽ��Q7��-a�;h��S������<�������;�����=������Q���6h���-a�X7���x   x   �7��Q���9�z��֧�6X��IX��֧�g���9�Q���7��fX���)�Q5T��|��h���Ǧ�G���6*��)�ž*�ž6*��F����Ǧ��h���|�I5T���)�fX�x   x   ���߭i�L��=׼t�� ���t���<׼M��ܭi�����7潾j��A��{m�h,��퟾񽰾3���I�ž�NȾI�ž4���𽰾퟾i,���{m��A��j��7�x   x   􌽕gC�a��j���ܔ��ܔ��j��a��gC�􌽫 Ž-��J�+��V�񂀾m���+���䵾�>��n�žn�ž�>���䵾+��h���킀��V�O�+�+��� Žx   x   g�o��W�ݼ��Fm����2�ݼi��)g��b��m~߽}I�'�:�Ymd�6���L���-����嵾l����-��n����嵾)���M���?���Umd��:�|I�r~߽�b��x   x   �;8�����8I��n��q��EI������;8��f���K���X�����|�D��k�̈�C���#-��"����������� ���'-��D���̈��k���D�����X��~K���f��x   x   JE��ɼЊ��1j�������ɼGE��M�F��ý=� �\c#���G���k�����> ��񟾽̦��"���̦��< ��������k���G�Yc#�7� ��ýK��M�x   x   ^3ڼ?[��%��%��_[��X3ڼ���G\�3��y+˽�%��d#�<�D��qd�O����0��2n����������3n���0��K����qd�>�D��d#��%��+˽5���G\���x   x   u�WQz���`�Qz�k򣼽~�W�#��Fd��ǚ�-˽� �,��[�:� V��m����o���]��o�����!�m� V�V�:�0��� �-˽�ǚ��Fd�l�#��~�x   x   1�v���J���J�L�v��맼��3f&�:Hd�u��y Ľ;`���N���+�n�A��@T�;a���g���g�;a��@T�i�A���+��N�5`��w Ľ��KHd�*f&���맼x   x   ��>�ر,�[�>�s>u�R[����#��L\�����]R��r�߽����s�f�)��7���?��B���?�7�o�)�}s����t�߽cR�������L\���#�"�s[��m>u�x   x   ����'�:�S>u��짼���S���#M��l���k���Ž0G��a���1������1���a�3G潏Ž�k���l���#M�X������짼*>u��:�x   x   .��T�����&'@��g}�_O��?ڼ�I�/�-�SS�=�y��N������p���w봽�ŷ�~봽p��������N��A�y�FS��-��I�LڼUO���g}�
'@�2��i��x   x   M��}�7��u�B�Ct��h���'¼�����/�.�L�J�)Ee�8�{��օ�Y��T���օ�9�{�-Ee�;�J�+�.������'¼�h��Ct���B���M����x   x   u��T��D4/���G��oj�e�������ȼq��+o
�5��/�1�<�2�E���H�8�E�>�<�/�4��>o
�[���ȼ����e����oj�i�G�F4/����H�����x   x   >@�E�B�g�G�x�Q��Fb��z����������}wм��I|�������	���	����<|����mwм~���������z�yFb���Q�U�G�"�B�c@�j3?�o3?�x   x   �F}�3't�[[j��;b��^���_��i�C�x��*���8��t����Ш��V��򟱼�V���Ш������8���*��>�x��i���_��^�`;b�s[j��'t�eF}��Ӂ�0����Ӂ�x   x   �7���S������r�y���_��K�t�>�f9�fW9�)�=�YC�ãH�}�K�`�K��H�.YC�߉=�qW9��9�n�>�B�K���_���y������S���7���ϰ������ϰ�x   x   ��ټ�
¼���|��j�h�r�>�;����u��Uϻ,�»<+��E��Q+����»-Vϻv廈�B�W�>�U�h�����
¼��ټ��CS��c���XS����x   x   �4�@��{�ȼ������x��8���S��Jk�����ӹ�d/���/��	Թ�5���Ik�|S�����8���x�������ȼ5���4��(��&���,���,��&��(�x   x   I�-���d����������59��L�%k�������7:���:�;���:�7:	���q$k��L��59��������B����C�-���E�ܸX���d�6i���d�ϸX���E�x   x   ��R� �.�&X
�&Rм���!`=��ϻ�z��M8:�*+;�Jh;_Jh;�*+;zP8:�{��ϻ`=����RмBX
���.�t�R���t�Ч������ek��lk������ͧ����t�x   x   �oy�l�J�5������۞��(C�sH»%�����:_h;yׇ;�^h;���:L$���G»�(C��۞����(��]�J��oy��/��=���ն������bĽ�����ն�A���/��x   x   T;��g#e���.��N������<oH�x໻�f���E;<kh;{kh;�F;cg���໻goH������N����.�i#e�^;������ƽH=ܽt5�L���R���s5�;=ܽ"ƽ����x   x   L����a{���<�,��\2��H�K����R\���:iQ+;��:�\��#���A�K�>2��/����<��a{�H����`½h�㽩w �����<����<�����w �[���`½x   x   1����ą�q�E��	��{��ۈK��޻�7����8:y�8:�� ߻���K��{���	�{�E��ą�/���4Kսr����.�?� ��{+��51��51��{+�E� ��.�p���4Kսx   x   dִ����٧H���	�?4��;qH�=D»�]��>���^�&D»EqH�"4����	�̧H����dִ�3�����n��Y2��^A�S�J��%N�_�J��^A��Y2�t����+��x   x   ʱ��n���E�������;+C��ϻ��j���j��ϻ(+C�"�������E�q��ұ����g?���(�@%@��VS��a��h��h��a��VS�>%@���(�o?���x   x   �ش�Sǅ���<�TV��t���$b=��A�?5��SA�Ub=�m���NV���<�Xǅ��ش�Q�vr�(.�`�H��`��r��P}�Ɩ���P}��r��`�c�H�%.�nr�X�x   x   �����i{�z�.���#!��79�������69�!���缆�.��i{��������:A�>.���K���f���|�'��z1��}1��'����|���f���K�B.�<A����x   x   �����-e����K\м���0�8�'��8����R\м���-e�����Rսc���(���H��f�f.����j9��V��c9����l.���f���H��(�b��Rսx   x   �B����J�p`
�����x���>���>���x����y`
���J��B���i½2���r�*@��`���|����"H��2���5���%H�������|��`�*@�o�@����i½x   x   �y��.�f�������h�j�K���h����Z��ݲ.��y��ʫ�!��5�C`2�+]S��r��)��;������������ ;���)���r�,]S�G`2�	5��㽟ʫ�x   x   zS����%�ȼ&����_���_���G�ȼ���vS�:���+ƽ �`� �*gA�'
a��X}��4���X�� ��������X���4���X}�
a�%gA�d� � ��+ƽ:��x   x   U�-�1��ϡ��R
z�^�_
z�������`�-�C�t�6+���Lܽ���S�+�n�J��&h�s����5���<���J���<���5��m����&h�{�J�P�+�����Lܽ2+��K�t�x   x   WB��¼3����Cb��Cb�F���¼VB���E�/���嶽�G�SG��@1�O1N�(h��[}�,��G��B�� ,���[}�(h�F1N��@1�VG��G�$嶽0�����E�x   x   :ڼ�b�� lj���Q�lj��b��@ڼL9�@�X�@��]�����������A1�.�J��a��r���|�73����|��r��a�/�J��A1��������X���<��9�X�P9�x   x   �J��?t���G���G�b?t��J���#�M�&�^e�r{��QvĽʬ��kI�Ո+�YlA�"dS�v#`�\�f�_�f�w#`�dS�UlA�و+�jI�����VvĽv{��le�L�&��#�x   x   8d}�M�B��</��B�d}�G氼�r����,��8i��|��1����L콿���� ��g2��2@�q�H���K�h�H��2@��g2�� �����L�8����|���8i���,��r��H氼x   x   �'@�M������'@��䁼�������0�,��e�����궽�Tܽ�� �3<�?�i�(��.��.�q�(�5�,<��� ��Tܽ�궽����e�8�,���������䁼x   x   ���T!�9���J?�'
������v���&���X�`����2��/6ƽM��x��� ��4L�t~�-L� ������T��&6ƽ�2��e�����X��&�jv�����+
���J?�x   x   ���h������J?�u偼R鰼�*�*?���E�j�t�C��:֫��w½.cս&�&�&�&�,cս�w½7֫�C��v�t���E� ?��*�d鰼~偼�J?�O��x   x   ����>�û�j������@�ھ{�잢�eμ�R��[��5�73P���g�(z�-����
��)���*z���g�A3P��5�[��R��[μ잢��{�o�@�؆��k�T�ûx   x   ��ûԻ�������9���g�GI��m����׼���ٕ��O&��*6�´A���G���G���A��*6��O&�ԕ�����׼����^I��r�g��9�>��4����Ի�ûx   x   �Y�d������0�U�0��|P�\�w��Z��7����Jɼ��伖4��Ko����������`o��4������Jɼ9����Z���w��|P�w�0�0����ݚ���Y�'�x   x   rw���P)�J��8))��9�.O��j�4e���y��������5��l�żq�ż5����������y��.e���j�GO�+9�C))�>��;)�����w�����x   x   k@���8�4�0�!)��k$��$�z)�@3��+A�>�Q�(�a��co�tx���{�4tx��co�M�a�n�Q��+A�;3�q)��$��k$�� )�f�0�4�8��j@��E��mG���E�x   x   ��{��xg�dP��9��$��a���+��� ����h��H	��4�T4��H	���H���� �L+����a��$��9�dP�Dxg�ԛ{�C��<��4<��C��x   x   )���&4���w�$�N�h�(���^�ڻFβ�b���;Ƀ�.�p���d�Xa�I�d�}�p�YɃ����β���ڻ��`�(��N���w�P4��7���?��#x������x��J��x   x   ��ͼ)����C���j�2�2����5�c�ʮ�1�p��z��t��83��8�|��Ѯp�`����c�����W�2���j��C��+�����ͼ��弒m���J �xJ ��m�����x   x   D-����ּ�x��N��|A��� ��e�����'���:��;�;��;��:��'�ؒ�Pf���� �(A�N���x���ּ+-��	��z�� �(�0�+�4�(�o����x   x   �D����)ɼt^���]Q����'���w�o���:�39;�h;R�h;�39;��:i�o����a���]Q��^��@)ɼ�����D�w/3�;6H��yW��_�ׂ_��yW�J6H�o/3�x   x   ��5�o��m������a�o���op���|���;[�h;ֆ�;@�h;j�;��|�uop�x���a������m�k���5�B�V�g�s��r���ڌ�Gi���ڌ��r��i�s�8�V�x   x   P�77&����l���/o��!	���d�/�8;��h;�h;#;��84�d��!	��/o��l�����B7&�P�s�y��$���V������0���0�����V��%����y�x   x   ��g��6��Y�~��@>x�2�Z�`����85�;�Q9;��;ө�8��`���=x�����Y��6���g����#_���к��˽�bֽ�ڽ�bֽ�˽�к�_�����x   x   Y�y�z�A���ݷż7n{�]��d�|�KU�:�W�:��{�%�d����n{�Էż���v�A�_�y��������ӽ�齅����$��$�����齛ӽ������x   x   �ŰG�����żAx��"	�Vhp�ˊo�a����o��hp��"	��@x��ż���ΰG��u����ƽ�-����5�V����Y�5�����-罧�ƽu��x   x   ����"�G�Ʋ�����4o���9���*p�Rp� �������4o���ϲ��G�����5���Q�Ͻ������O���$���)���)���$��O������[�Ͻ6���x   x   ����8�A�X]�r����a�\��]��w�c��\�����X�a�
r��D]�6�A�����L���Lӽ!��)v���#��A1��9�D�<��9��A1���#�0v�!��AӽJ���x   x   �z��6����p���dQ��� �ү������� ��dQ�u�����6��z�Ex����Ͻ�"�����`�(��J9�?E�G8K�J8K�CE��J9�[�(�����"���ϽHx��x   x   ��g��>&��x伬e���A�����ڻ���A��e���x优>&���g�	�����ƽ�����w�k�(��
<���J��_T�"�W��_T���J��
<�k�(� x�������ƽ���x   x   �!P�����4ɼU��h�2�J����2�U���4ɼ����!P�������5�	���#��L9���J��W�p^�u^��W���J��L9���#�	�%5�������x   x   �5����������j���(�4\���(���j���������5���y��g���ӽ����T��E1��E�wbT��^�Oa��^�zbT��E��E1��T�����ӽ�g����y�x   x   /P�Z׼N���O��$��$��O�*N��i׼*P�,�V�-.���ۺ�Ǥ�o�"�$���9�I=K��W�0^�,^��W�L=K���9�!�$�p�ä齉ۺ�4.��(�V�x   x   �B��1�����w��9��j$��9���w�����B��>3� �s��a���˽������g�)�Q�<��>K�eT��W�&eT��>K�M�<�g�)��������˽�a����s�>3�x   x   Lμ;A���rP��&)��&)�sP�NA��Iμ����GH��}������qֽ"-�H����)�9�9��E��J��J��E�;�9���)�I��#-��qֽ����}���GH����x   x   ����Y�g�"�0�ʍ�1�0���g�����漎����W�z猽�?���$ڽ	.��!�m�$��J1��R9��<��R9��J1�l�$��!�.��$ڽ�?��}猽s�W������x   x   ��{�G 9�2�2�� 9���{��,��r���n�(���_�Bw���@���tֽ���J��Y�"�#�%�(�*�(�!�#��Y�L�����tֽ�@��Bw���_�|�(�|����,��x   x   À@�4��ى������@�zS��3����Y �&�+���_��錽����˽���������q������������˽����錽��_�+�+��Y ����~S��x   x   8��׫������z���E�>N��~ν��Z ��(�f�W�􁅽�g���㺽|ӽB�����3���3������B�tӽ�㺽�g������c�W��(��Z ��ν�>N��#�E�x   x   Eo�+Ի=n�K���G�)O��ב��	���o���OH��s��5��2q�����ϱƽ�Ͻ�*ӽ�Ͻñƽ���>q���5����s��OH�q�����ő��O��n�G�M�x   x   ��û,�û�%�7�k�E��U���1����H���G3�B�V���y�S%��y��������������������G%����y�H�V��G3�P��w漣1���U����E�7�%�x   x   �d���9��t᲻�߻>$�� :���m��:���~���ܼ�7�-v�g�#�Tf0�w�8��i;�f�8�Yf0�k�#�/v��7��ܼ�~���:����m�� :�$���߻ⲻ�9��x   x   �4��r��F��Rử�	�_p*���Q��!�����G���
RѼ�&�8� ��{�P��g���{�'� ��&�	RѼI�������!����Q�Op*���	�������5��x   x   ղ�����?̻{c�E���V��43�s%S�w�����P���D���׿��ȼ�˼��ȼ�׿��D��{P������w��%S�V43�XV�l��ec仞?̻+��ղ�8կ�x   x   n�߻�ởY�b�����
����m_&���;�w�R�N�i�e`}���������E`}�$�i���R���;�n_&���]������a뻛Y���k�߻Ҩ߻�߻x   x   ����	�S��,������<5껉���A��aR�J��)����#�g�)���+�y�)���#�N��u��=R��A��o���4�A��#���{����	�e�YF���9F�x   x   !:�$Z*��D����b(�5�λ��ݎ����ƥ��!����4���b��jb���4��[���R������%�������λt(�����D��Y*�Q:��E��K���K��E�x   x   p�m�>�Q�53�J	�m��-��l����c���5�������,񺽘��-�����L�5��c�+������M��C	��3���Q���m��ف�"T`��%�ف�x   x   -%����:S��D&�����u��hc�� ���S�ȭ�7J�:��T:��T:D�:F��7<�S�l� �hc�[v�����D&�hS���	%����������ɺ��ɺ��������x   x   d�����v�t�;��8���5��ZS��4:d��:�;';Ԯ;���:�4:�ZS�֡5��𪻙8���;���v���d��Z�ѼP�ܣ�=����P�7�Ѽx   x   haܼ.���w�� �R�����x���r�7��7M��:��:;],_;F,_;��:;���:Ѻ�7�q�|x��պ�!�R�$w��+���laܼ+2 ��^�^d�\5 �A5 �Ld��^�(2 �x   x   �%�D2Ѽ�5��bi�Uo�ǋ�����M�:��;8_;{6v;�7_;��;��:���؋��9o�
bi�k5��J2Ѽ�%�����-��>�εH�p]L��H��>���-���x   x   Ub���E'���0}��#�����އ��U:E'';|?_;?_;�'';0�U:%������0�#��0}�^'����Ob��	1��qL�wvc�:t�!�|��|�9t�tvc��qL��	1�x   x   N�#��p ���������)��'����麣�U:��;��:;�;!�U:/��a'��?�)�:�������p �M�#��sG�Z�i��!����������R���������"��X�i��sG�x   x   �P0�i��ȼ�Չ��+��'��m����:���:� �:&�:����'��y�+��Չ���ȼi��P0�k<Z�rၽ���*��f����������k��������vၽi<Z�x   x   �8����˼�։�Y�)�����a����7+�4:���7�������)��։��˼����8���g����Z���_���Eǽ�iѽ��Խ�iѽ�Eǽ�_��Y�������g�x   x   U;���s�ȼ��D�#�����Oh�j�R���R��g�k���z�#��򅼃�ȼ���T;�5�n��y��+.��2�Ž�$ڽ���T��U���轍$ڽ-�Ž+.���y��.�n�x   x   :�8��k�꽿��7}��s�y��U�5��e �[�5��y���s��7}�ݽ���k�H�8���n�Ȳ��w����ν��罦
����?��
���
�������νw��ʲ����n�x   x    U0��t ��-���ji�Y��f��Qc��Qc��t��ki��-���t �#U0��g��{��7x���ѽ��KL� ��ZN�WN����PL����ѽ1x���{���g�x   x   v�#��=����R��<��r��s��Hs���<���R�=���q�#�GCZ�`��o1����ν��G���1���O�5�����G����νl1��V��MCZ�x   x   �i��=Ѽ!�� �;�%!��������Q!���;�*���=Ѽ�i��|G�W恽z��+�Ž���M���>��������=����M�߬�&�Ž���X恽�|G�x   x   �-�䑵���v�TM&����ڭλ���IM&���v�ߑ���-�g1��i�D	���f��l+ڽ��������� ��h �� ���������k+ڽ�f��D	���i�f1�x   x   Kqܼ�����S�4�M(껝(�*��S����Bqܼ`���~L�u)��}���NǽX��.���Q��R������R��Q�,��b�轠Nǽu��r)���~L�^��x   x   s��l��['3� ��x�����V'3�_��s��J< �z�-�#�c����x���~tѽ��W���R����@����R�]�� ��mtѽz�������c�v�-�L< �x   x   �2����Q��N���������N���Q��2��.�Ѽk�G/>��+t�R�������8�Խ�����a��n�o�c�������C�Խ����J����+t�O/>�k�-�Ѽx   x    �m�2i*�w���e�x���h*�#�m�����f漿r�{�H��|��^��󥶽Twѽ�车��LR��L�JR������Qwѽ���^���|���H��r��f漊��x   x   �:���	��e仞e���	��:�聼w��~��vE ��pL���|�t���7��� Tǽ�2ڽB�罳���<���2ڽ$Tǽ4���v�����|��pL�iE ����x��聼x   x   �!���H̻(��!�w�E������ߺ�Y���F ���H�1t����G��`n����Ž��ν��ѽ��ν��ŽWn��J�����1t���H��F �+Y���ߺ�y���~�E�x   x   �߻\#���#��N�߻KX���K�r��Ẽ~��=v��4>���c�8/������!��D<������z���A<���!�����0/���c�
5>�Gv�]���ຼBr����K�YX�x   x   �䲻���䲻�߻7��B�K��������m漠p�`�-�a�L���i��U�����>���&���M�����i�k�L�^�-��p��m漥��{���K�A���߻x   x   P<���<��&䯻6�߻]Y�!�E��끼���ѼIC ����r1�_�G��TZ�/�g���n���n�3�g��TZ�Y�G�q1����MC ��Ѽ���끼3�E��Y��߻�㯻x   x   ��`�� m�`a��$稻�gջ�y���*��S�-뀼`ə�x2����˼W%Ἲ �N���f^ �?���� �[%���˼q2��hə�)뀼��S���*�z��gջ�樻�a��� m�x   x   �m���}��o��T����˻������4��^W��>|�Ꙑ��ӡ��h��7����������D���h���ӡ�Ꙑ��>|��^W��4���ӏ��k˻˹���o����}��m�x   x   �X���j����z��ͩ���dڻDR������=+�bD�OA]���s����Ո�7⊼�Ո����s�oA]�
bD��=+�����Q��CdڻO���z��i��j���X��._��x   x   ר�����s���5���f�� �����λ�,��6 �(������*�+�4�m�9�|�9�T�4���*������6 ��,廦�λZ����f��.5��Ds��<����֨��$��)%��x   x   �Nջ��ʻW���|^������֢��j��`��d y��t�ʻK�ֻr�޻�H�6�޻A�ֻ��ʻy��g
`��mj��֢�c����^������x�ʻ�NջI,ܻ��޻,ܻx   x   �g��p��^Kڻd|��	͢��c��bw��a���U�4�R�QT���W��Y�R�Y���W�5T��R���U�Ma�cw��c���̢��|��JKڻ^p��"h�uN�����YN�x   x   �w*�����.��8hλ%X��8�v�*�6�ѕ��ῺZ@��|`Y��q5�N*��r5��`Y�G@��nῺ��f�6���v�#X��4hλ.������w*�\;���E�wDI���E��;�x   x   ��S���4�7|��kD���`�����Gh�}_9�ӏ#:!��:��: �:ղ�:s�#:�|9�Gh���?�`�RD���_|�Ù4�;�S�7�m��X��-X��%X���X��5�m�x   x   �؀�a=W�!+�{ �Mʰ�[�U�#���E�*�㨐:o��:�];[~$;];0��:Y��:�*������U�fʰ�� �� +�F=W��؀����1����*���z���*��<���󮓼x   x   ����u|��@D����M��ԌR�j茺��#:���:�2; N;6 N;��2;���:�#:�猺�R��M��]��@D��|�����\?����ȼ�Iؼ�|�o|༛Iؼ��ȼX?��x   x   ���郐��]����4�ʻ�4T�H�X�M��:r;�N;P2_;�N;�q;���:��X��4T��ʻ����]�냐�����1Լ�m�6�7��\�M��6��m��1Լx   x   �w˼���B�s��*�^ֻ�AW�J�4��i�:G�$;�N;FN;^�$;�j�:׃4��AW�%^ֻ�*�U�s�����w˼���[��C���(��.���.���(��C�[�ն��x   x   qἌO���܂�m�4�YJ޻�`Y��)�0p�:�y;��2;�y;p�:�)�b`Y�J޻��4��܂�yO�����P	�y!�U�5�GOF���P�cT���P�EOF�V�5��!��P	�x   x   �������9��haY��{4��	�:U��:���:	�:ez4��`Y�gỚ�9�w�������eM2�j�L�
wb��Ir�P�z�k�z��Ir��vb�g�L�bM2����x   x   ��������X͊���9�oL޻�BW�swX��0$:�ܐ:�0$:VwX�.CW�nL޻��9�c͊���������}�� �?�;a_�0{����vv��Gۑ�gv�����(0{�0a_�"�?����x   x   CP �ƍ��+�П4�Sbֻ�5T��׌�`��(���֌��5T�kbֻǟ4�+�����<P ���#�9uH���l�3C���K���f�����������f���K��6C����l�&uH���#�x   x   ����)��߂���*�ةʻ�R������g�����H�R���ʻ��*��߂�%�������#�mK�)t��l��a}���ث�h\���H��k\���ث�_}���l��0t�2mK���#�x   x   		��T���s����XS���U�bs�2s�b�U�gS������s��T��
	�g���wH��t�&���#L���ĳ�9�����Ž��Ž2����ĳ�)L��$����t��wH�l��x   x   ���¡��%]���4ϰ�L�`�֌6���`�Kϰ����%]��¡���K����?���l��n��(M���}���yŽ1Ͻ�Gҽ>Ͻ�yŽu}��+M���n����l���?�K��x   x   ��˼���$KD��% ��G����v���v��G���% �8KD�����t�˼�V	��S2�h_��F��Y����Ƴ��zŽ�,ҽ��ؽ��ؽ�,ҽ�zŽ�Ƴ�U����F��h_��S2��V	�x   x   /$��>'|�e++���)Y���[��IY����Z++�<'|�1$��%���N!�5�L�u9{��P��9ݫ�ڝ���Ͻ9�ؽ�*ܽ9�ؽ�Ͻ۝��7ݫ��P��t9{�=�L�R!����x   x   3���vLW�̅��pλ�ˢ��ˢ��pλׅ�mLW�1����?Լ�c�W�5�@�b�����l��b����Ž�Kҽ��ؽ��ؽ�Kҽ��Žb���l�����:�b�S�5��c��?Լx   x   �‼��4��>��Ƃ��9~������c>����4��‼�L�� �HN�[F�Wr��}�������O����Ž�Ͻ�0ҽ�Ͻ��ŽP�������}��Wr��[F�JN�'��L��x   x   ��S���RXڻ"b��:b���Xڻ޳���S�λ��7�ȼw@��(���P��z��㑽"����d�������Ž�Ž�����d������㑽(�z���P���(�v@�.�ȼѻ��x   x   ��*�Ƅ��!���7��社�����ч*��m�n���]ؼ!���.�sT��z�����o���᫽ͳ������̳��᫽�o������z�
sT��.�(�� ]ؼu�����m�x   x   �u��˻�z��{���˻�u�;�?f��$<��h�༅&�R�.���P�E\r�Љ���U��ʆ���T���T��ǆ���U��ω��;\r���P�a�.�|&�X��&<��>f��;�x   x   $dջ��������ƹ��#dջ�^�B�E�3g���������N����(�-aF�5�b�D{�M��3v������>v��M���C{�:�b�5aF���(�@����ō��(g��A�E��^�x   x   �樻�s���s���樻[Eܻ"�']I�:h��?��bؼbD�T�<�5�c�L��t_��m�|t�lt��m��t_�n�L�7�5�T�sD�(bؼ�>��6h��M]I��TEܻx   x   bc��x�}�Qc���6����޻)�U�E�+i������)�ȼ(���j��!�z_2�y�?��H�/~K�(�H�}�?�s_2��!��j�1���ȼ����Ni��?�E����޻�6��x   x   $m�$m��i���6��Gܻ^a��;���m����V���LԼ�����`	�e��:��ś#�ƛ#�5��`���`	������LԼ�V������m��;�ya�DGܻ�6���i��x   x   ��1�Me:���S��h~�gʜ��»�X������0� Q�-�q�P���U{��BT��W?��
���g?��DT��V{��T��� �q�Q���0�����X�`�»-ʜ��h~���S�Ke:�x   x   m`:�.:E��	[�6�{���������ąѻ,������p*�:!B�4X�3�j��kx����U��pkx�K�j�4X�A!B��p*�����+���ѻ9���������{�!
[�S:E�K`:�x   x   ��S��[�:hg���y��B���홻4D���(ɻ�滑6����rE!��,��U4�t�6��U4��,�lE!�����6����(ɻ&D���홻uC����y�egg�r[���S���Q�x   x   �R~��{�	�y�Py�[�|��v���[��]*��B7��s>��vqͻ��ݻg)������N)���ݻ�qͻc>��57��R*���[���v��,�|��
y�[�y���{��R~�������x   x   .���h瓻M8����|���i���\�!~V��W�,`��@m��c|�)/������΋����Z/���c|��@m�z,`�>�W�~V�ߤ\���i���|��8��瓻����v��_u���u��x   x   �w»!���<ܙ�jj��,�\��)8�Mp��;��������n�0�麋!�7"���Yn�|��'��Q;�Hp��)8�\��j��1ܙ�򝯻�w»�?л�y׻�y׻u?лx   x   8�hѻ�+���H���dV��c���Ӻ/B�����S���}�� X8I��8lX8р���S��r��VB����Ӻ�c�"eV��H���+���hѻP8�d��K�5��K��d�x   x   *������ɻ�����W�H#��*��l�/��i�9G�|:�:��:$�:��:��|:�i�9��/��*���"���W�����ɻ�����ʯ%��k3��:��:��k3�ί%�x   x   ��0�������D�_�����]{����9��:��:5";�;%";&��:���:z��9?z�;����_���ٛ�ӵ���0��tK��v`�y�m���r���m��v`��tK�x   x   �Q�^V*�������m�+��}\����|:��:+�#;��7;��7;C�#;��:{�|:�]�����Tm�C����xV*��Q���t��-���쓼����m����쓼�-����t�x   x   ��q��B�D���Fͻ�|���ߝw��>�:�0;�7;�CD;�7;�0;�>�:Чw�r� |�Gͻc��lB���q���������=J���B��̮���B��J��򣣼����x   x   ����X��)!��ݻi
���?�(�b8EK�:��;�7;�7;��;�K�:p�b8�?�f
����ݻ�)!��X�"���.���PU���Ӽ�)��8��8��)�*�ӼNU��"���x   x   h��b�j�M�,�����ꉻ}�꺬z�8�O�:�6;»#;�6;�O�:u�8ӫ�뉻���e�,�]�j�h��zط���׼Ӕ�+��������(����󼺦׼�ط�x   x   �@��0Ix��84���ר�����c8,K�:�!�:�!�:4K�:�c8<�꺓������84�4Ix��@����Ǽ���Y����)g!�h�&�m�&�&g!�����Y�����Ǽx   x   �+���k�%�6�y��6쉻q@�#�v�}}:��:�}:�v�t@�z쉻���6�6��k��+���[Ӽ�.��)}���&��K5�u�>�ӪA�p�>��K5���&�}��.�� \Ӽx   x   /���m�;4����8����\'��� :� :(����������:4�&m�@����aټ��7�b^3�c�E�W;S��8Z��8Z�[;S�^�E�p^3��7����aټx   x   �-���Mx�V�,�=�ݻ&|�ъ��Q��.�5R�v�꺄&|�1�ݻ{�,��Mx��-���bټ����!��U;� �Q��sc���n�*�r���n��sc� �Q��U;���!���bټx   x   SD��Z�j�R/!�vNͻ�
m�u��������������
m��Nͻ:/!�>�j�RD���_Ӽ� ���!�>��X���m�p}�aЂ�cЂ�p}���m��X�">���!�� ��_Ӽx   x   Um��vX����J ����_�R���ӺX���_� ������X�Xm��Z�Ǽ�4���:��W;�AX��Zq������∽0���∽ߒ���Zq�BX��W;��:��4��K�Ǽx   x   h���JB�f&�a����W��Y��Y���W�z��p&�,B�i����߷�&�����b3���Q���m�����[��� ^�� ^��^���������m���Q��b3������෼x   x   y�q��`*� �����dV�88�ydV�����滊`*�|�q�����°׼G_���&�s�E��yc��t}��䈽
_��Θ��
_���䈽�t}��yc�p�E���&�Q_�Ȱ׼����x   x   jQ�����ɻ�M����\���\��M���ɻ����Q�����V`���������S5�/CS��n��ӂ�����_���_������ӂ��n�0CS��S5�������U`������x   x   ��0�����5��rm��#�i��m���5�������0�{�t�8�����Ӽ���o!�܉>��BZ�`�r��Ԃ�^戽���Y戽�Ԃ�[�r��BZ��>��o!�����Ӽ-���v�t�x   x   ��KxѻQ䙻��|��|�I䙻(xѻ��?�K��8���W��:�0����&���A� DZ�N�n��y}�!���'����y}�T�n�DZ���A���&�5�� :㼳W���8��;�K�x   x   WM𻴪���>��`y��>������FM�ʾ%��`�����dR��<K�4#���&�w�>��GS��c���m�dq���m��c��GS���>���&�+#�<K�_R�������`���%�x   x   ��»��0�y���y���s�»�q�|}3�wn�ӝ������L�.��[s!��X5�0�E�`�Q�eX�`X�g�Q�2�E��X5�Ys!�2���L����ʝ��Nn��}3��q�x   x   (ǜ��{��mg��{�'ǜ�.Uл�Z��:�M�r��LU���>����L����&�gk3�	b;��>�
b;�ak3���&�J������>�4U������r�r��:��Z�Uлx   x   h~�Q[�[� h~���׻����:�dn����]����Ӽ+��f�݉��D���!���!��D�׉�f�4���Ӽ]�����&n���:���7�׻醢�x   x   ��S�;AE���S�������ȓ׻�\�Ӂ3�;�`��=������Gj��m�׼{���F���*�7��*�G��{��g�׼Hj�������=��Q�`��3��\���׻������x   x   �g:�xg:�T�Q�A��m���kYл#v���%�9�K�4�t����� ������ǼrӼwټwټrӼs�Ǽ����������>�t�E�K���%��u��Yл����k��m�Q�x   x   i����J%��]@���e��I������B�ǻ)��/8
�h_�Ǖ1�	sB���O�q�W�3�Z���W���O�sB�ٕ1�a_�8
����S�ǻ֠���I��J�e�h]@�kI%����x   x   ����r��(��I<�LuV��w�i���맻��»�g߻	#�� q�~��J��4"#��!#�#�����!q�#���g߻��»�맻O��f�w�QuV�>J<�0�(��s�c��x   x   �A%��(��h.��67��D��U�'�m�ޛ��r��V��j���#ͻ��ڻ���V��D���ڻ� ͻD����V����͛����m�k�U�D��67��h.�(��A%�9/$�x   x   �N@�^><�@07���2��0�
3��:��3F�^�V��rj���~�Bш���I�������Jш�j�~��rj���V��3F��:�9	3�,�0�_�2�[07��><�jN@�0�B�ȅB�x   x   ��e��aV�l�C�]�0���L��֍����+����
�v�����t�st �Uu�G�����
����м���������9�0���C�aV���e��[o�۷r�r[o�x   x   ^9��Amw���U���2�ܗ�2�*��������v�G[���N�K K�H�J��J���J��N��[���v�垓�����/躣����2���U��mw��9��(蔻<�������4蔻x   x   �������`�m�y�9��|����zIW�� ���>o���~93(�9%:H�:)&:�%�9��~9��m�+!���JW�󰷺}���9��m��������S���t>ĻKȻ>Ļ{���x   x   �ǻ9ӧ�����dF���g~���๹�׏9�-G:竑:���:ע�::)��:ج�:4.G:�ԏ9๹}�����rF�V���Jӧ�0�ǻC`���� �) �;���@`�x   x   :�컫�»q���R�V�����tv��f2�7JG:AͰ:���:94;G�	;�4;��:̰:EJG:Wv0�wv�P���V�������»@�컡���W�>� ���#�3� ��W����x   x   �$
��D߻�8��=@j�X�
���Z�(�9�ő:[��:y�;��;��;��;G��:Ǒ:-�9וZ�y�
�/@j��8���D߻�$
��g"���6�E���L���L�-E���6��g"�x   x   �I�����ջ��~�����N���9��:{>;L�;l�';S�;?;k�:V��9�N���J�~��ջ������I���<���W��fl�b�y�4*~�~�y��fl���W���<�x   x   6~1�\���̻����9���eJ���:�˾:��	;�;R�;f�	;�ʾ:�:�cJ�A��Ȳ��7�̻$\�Z~1���V���x��j���,͙�͙�ބ���j��+�x���V�x   x   )ZB�p����ڻ\쏻fA�W�I��N	:�;:�C;�;�C;�;:�P	:��I�WB��돻H�ڻ���ZB�aOn���9$��MW���b���~��c��KW��$���󋼄On�x   x   8�O������㻉䓻A �=�I��:;�:տ�:u��:��:d�:��I�*@ �r䓻������-�O�J�l���f ����¼Taм�p׼�p׼?aм�¼� ��_���;�x   x   �W�)#���� 哻�C�dJ�M�9_֑:|�:�֑:��9lcJ�D�N哻;���#�&�W�C���,=�����A�ּ_�������������\��ּ���A=��=���x   x   ��Z��#����P���\
N�?�9�wG:WwG:=�9
N�"��nA���#���Z�Ҥ��a��#�ɼ4漍���>J�k��l��@J�����K�)�ɼX��㤋�x   x   ��W�k���ڻ`���t����Z�0��NM�9�����Z�N��e���.�ڻ�����W������X���pϼ����2�r^���:����p^��2�v�＄pϼ�X������x   x   ƉO�����̻9�~���
��fv�C���]���Mhv�R�
�ٶ~���̻���ƉO�����R���qϼ�B�
����H�!�%�&�7�&�X�!����
��B��qϼ/������x   x   �`B�Wa�ݻ�#Ij����~q��>W��p�����Hj�uݻ�ja�t`B������@����ɼ[���
���&�Uw.��41�<w.�&�	��
�'�Ｚ�ɼ�@������x   x   ��1����@���V�����ɟ��h�� �V��@������1��Xn�����c����+5�����&�1���6���6�1��&����<5���A�������Xn�x   x   $R�Q߻V����F�jz�"躘z��F�Y���(Q߻(R��V�����g'����ּ����a�B�!��y.���6�1n9���6�sy.�G�!��a������ּ|'��������V�x   x   Q-
���»e�����9��������9�7���z�»v-
���<���x�<,����¼�� O�[��L�&�81���6��6�81�X�&�a��O�����¼,����x��<�x   x   ���ݧ�k�m��2��y���2�f�m�ާ����s"���W�Os��$a��Llм����b�����w�&��{.��1��{.�r�&����k������;lм(a��gs��|�W�s"�x   x   �ǻO��*�U���0�{�0���U�&���ǻ��G�6��wl�����n��p}׼Q���T��W����!�e�&�f�&�{�!�k��]��.���n}׼�n�������wl�_�6���x   x   R���Q|w�H�C�3�2�r�C�3}w����"s⻆d�.E��y��ؙ�׋���~׼����Q��e���������e��Q�����~׼܋���ؙ�ٳy�E.E�zd�s�x   x   �D��XnV��47�57��mV�D����������г ���L��?~��ٙ�@q���pмb鼴����:�D
�F
��:�����e鼗pм)q���ٙ�@~���L��� ���������x   x   %�e�yH<��k.��H<���e������QĻ�& ���#�T�L�ȷy�2���f����¼~�ּ��2��qQ��；漠�ּ��¼f��@�����y�V�L� �#��& �QĻ����x   x   0\@�=�(�͚(�\@�xqo����`Ȼ( �f� ��2E��~l��x���2��O0���$��$�ɼ�ϼ�ϼ9�ɼ�$��90���2���x���~l��2E�8� ��' �Q`Ȼb����qo�x   x   cJ%��w��J%��B���r������TĻ���gi���6���W���x�"�������L��m��3g��S���L������7����x���W���6��i�.����TĻ�����r�7�B�x   x   G�����8$��B��so�Q�������|���f|"���<��V��jn�T ��f����������h��S ���jn���V�$�<�a|"�����|�ͥ��<���`to���B��8$�x   x   w��td�0��<���.(��HC�#�c���N-��Hݰ���ǻ��ݻ���������W$����������Ϧݻ�ǻ�ܰ��-����/�c�IC��.(�%�����gd�x   x   u`�3���k�O��rQ��-�pC��=]��z��A��3��$���x���o��ƻ�ƻ�o���x��.���2���A��J�z��<]�C��-��Q�a���k��4��X_�x   x   ����h���/
���� G�J���,��>��lQ��e��Dw�����ܭ��pL��&�������6Dw�le��lQ��>�e�,�K�hG�$��*
���<h�B��ڤ�x   x   ���҉���=o �Z0���A�j������2�
����B�Lq$�F`(��_(��p$��B�Y�f�
����x���j�;?��0��ho ���O��0��TF�?F�x   x   ) (��D�+��'&��R�ֺ2q��.���y���t��ɑ����J,������Y��I���O-��9��ȑ�?u����z����q��}�ֺ�%��2��%D�} (�'�0��q3�҉0�x   x   �3C�2-��7�$,�
f��ʘ��kfF�/���2����l�؁(����E��YA����e|(���l�64������eF�����2f���*��7��-��3C��S��U\�aV\�`�S�x   x   ��c�~C��4�WI𺚆���OF�Jգ�W�O8*��9�	:��+:�8>:�7D:9>:��+:��	:O��9�O8@ף�aQF�����QI��5��C���c�<�}�l��]���k��6�}�x   x   M℻4]��,�����㘺����Q8O|:p�d:2�:��:c�:��:��:�2�:F�d:{:6'Q8����㘺{���z�,��]�s℻8���Z)��F��?F���)��.���x   x   ����z�?�=�#��I��ֲ���ի9r�d:�.�:���:!�::��:�!�:#��:�-�:<�d:�ث9W����I�������=��z����xL����ƻ�qӻN�׻�qӻ��ƻ�L��x   x   /Ű��+��FQ��_
�N���h�k���	:nC�:���:���:�;;��:l��:�D�:��	:v�k�(����_
��EQ��+��Ű�!#ѻ����
���~��~��
����_#ѻx   x   ��ǻq��l�d�Z��䔺m'���+:v1�:/�:
;U5;
;
0�:<1�:��+:k
'�E䔺�����d�?���ǻ����T	�r��'l��\"�Hl�z���T	�c��x   x   Z�ݻ�뫻(w�x��뙺�����>:(�:e��:;;���:� �:�>:����뙺��pw��뫻��ݻ�����0�.�S�;�gB�gB�!�;�_�.�;�����x   x   ���]��r݂��H$�%T�������D:��:�5�:|�:q6�:��:܊D:9����U���G$��݂�2]��f��=g�>�.�"�E�I�W�fJc��3g��Jc�H�W���E��.�Ng�x   x   Gs���S������Z7(����������>:8�:��::�:�7�:�>:����_��7(������S��+s��-��R�>�x[��yr�V���������L��� zr��[�O�>���x   x   �s�ƻ�4���7(��V��:��.�+:�O�:A�:?P�:�+:���UW���7(��4���ƻ�s�ش'�?K�yl�ք�?:���z�������z��8:��ք��xl�ZK�δ'�x   x   ���ƻ3���CJ$�!��&��
:��d:��d:
:
�&�-dJ$�����ƻ�.�+���R�W�x�
����U��I���4(��:(��N����U�����W�x���R�E�+�x   x   Au�xV��6���+��唺Wlk�]�9��:g�9Pdk�s攺e�>����V��Au��+�+�U�:��⠓�m������~K���E��fK������n��ޠ��.���U�*�+�x   x   Px���a���w����[�������;S8�KS8z���9�������w��a��bx��x�'���R�����������5��w,Ƽ p̼p̼�,Ƽ�4�������������R���'�x   x   ��񫻄�d��c
�ZH�����H������H���c
���d��񫻬��O���K�jy���������м���˼-xռ,�ؼ
xռ��˼�м����n����y��K�F��x   x   6�ݻ!���NQ�T�������1F�4F�"���4��iNQ�� ��C�ݻ�l�X�>��l�2㍼@	��47��/�˼/�ؼU:߼c:߼D�ؼ-�˼%7��U	��5㍼ml�R�>��l�x   x   ��ǻ�2���>�R���/���녋����'����>��2����ǻ	����.��	[�}ڄ�:Z��֣�� 0Ƽ�zռ�;߼��⼲;߼�zռ	0Ƽӣ��4Z��vڄ��	[���.����x   x   �ΰ�|�z���,�dK�]���\��TK�z�,�R�z��ΰ����	����E�y�r��?�����	Q���t̼-�ؼ.=߼=߼4�ؼu̼Q������?��v�r�]�E������x   x   k"��X)]�j;�)𺑆ֺ*�};��)]�7"��0ѻ]	�7�.���W�ح��偗�L/���L��`v̼`}ռd�ؼn}ռWv̼�L��\/��恗�Э���W�P�.��\	�0ѻx   x   넻�C�i<��#���"���;�4C�넻�X����|��T�;�1Xc�J��� ��z0��lS���3Ƽh�˼l�˼�3Ƽ�S���0��� ��H��(Xc�G�;�o��I�뻑X��x   x   ��c��-����m ����w-���c�_����ǻ����w��tB�4Cg�$�����t¦�����@=���׼�:=������d¦�����7��JCg��tB��w����ǻc���x   x   AC��K������J��@C���}��6��F�ӻ����i"�6vB��[c������C���_�����ؚ��ݚ�����|_���C������g[c�?vB�j"�~���ӻ 7��L�}�x   x   *(���͛�z���*(�o�S��w���U����׻���kz�K�;�+�W�(�r��߄��鍼l���ᣕ�V����鍼�߄��r�M�W�p�;�Sz����>�׻�U���w����S�x   x   ���^l��k�.��j�0�8i\�j��1W����ӻ$��.����.���E��[���l��y�������y���l��[� F���.���5$����ӻW��j���i\���0�x   x   ��9�����P���3��k\��y��`;���ǻ��nc	������.���>�7$K� �R�̫U��R�"$K���>��.����c	��컏ǻz;���y��k\�&�3�OP�x   x   �e��d�Ԫ��P�g�0��S��~����Ub���<ѻ�����"x����Y�'�e�+�d�+�o�'����	x����s�ﻎ<ѻb��+���P~�ϬS���0��P�֪�x   x   ,ź�nȺ�"Һ��ẆR��h	��
��S-���B��Y��p��#��s���I��/Ř�c��"Ř���k����#��m�p�ƑY�H�B�T-�Z
�h	�
R�����#Һ�nȺx   x   �lȺ��ʺm�Ϻ+6׺S'�I�Ek�oV�+�=�*���9��G�w9S���[�|`��`�]�[��9S�ܖG�r�9��*�%��U�2k�MI�'�A6׺ӸϺ��ʺPkȺx   x   �Һ��Ϻ�X̺[ɺa'Ⱥ$�ɺ!]Ϻ{�غp庡���1j��	�&����V������-�	�Wj�W����p庺�غ�]Ϻ@�ɺ�&Ⱥ>[ɺPX̺�Ϻ�ҺR�Һx   x   V��
-׺�Uɺ�C��䫺�韺t�����ּ����������;)��A���c8��9��x���)��W���橕�ɼ��7��t���蟺w䫺�C���Uɺ�-׺�ậ�纜��x   x   �@���⺼Ⱥ�ݫ�4ᏺ��l��QA�+��7�Sp���V�߹U?߹x߹|=߹w�߹V�乥n� 7�	��eRA� �l��ᏺ�ݫ��Ⱥ��FA��ڛ���k��x   x   e[	�-2�P�ɺLܟ��l��F�����y�����7<9p~b9�܇9���9$��98އ9P�b9�69��7�������E���l�|۟�2�ɺ3�,[	�J���8��8����x   x   ����[��BϺ8_��?5A�덷���0���9R]:0�+:3�G:�W:P|\:��W:��G:r�+:�^:���9i�0�����5A�&_���CϺ{[�����,��8�ܛ<��8���,�x   x   ?-�2C���غ���������\��9�~ :�2f:VO�:�t�: L�:M�:|u�:'O�:h2f:Q~ :y��99���������غC�?-���F��[Y���b���b��[Y�-�F�x   x   �B���G���������7Pw:�>f:uڙ:��:F�:��:�D�:�:�ڙ:l>f:�w:���7T��Ù���G����_�B��Ld�DA~�S�� ��=S��CA~��Ld�x   x   AuY���*�C}�����f��	9�,:�Z�:�:�W�:a�:�:X�:��:�Z�:�,:9?�򹓁���|����*�&uY��́�1���l��֥��ե��l��#��3́�x   x   �kp��9��O�Yu��\乵lc9�*H:태:EO�:l�:�H�:g�:�N�:���:J*H:Glc9�[�.u���O��9�$lp�^ˑ�hꧻ�����û��ǻ��û��>ꧻ?ˑ�x   x   ���)wG���	�����tW߹:_�95�W:Q^�:���:�
�:;
�:���:_�:�W:�_�9�V߹<�����	�MwG�|���N��-����ӻ�#�_��i�뻍#㻊ӻH����N��x   x   ���.S����؄����޹��9ٱ\:�`�:*R�:�`�:OS�:�`�:��\:G�9��޹|������?S�����:`����ϻE���u
�	���E�`�ϻ`��x   x   U����y[�C��i����޹��9�W:���:%�:�$�:׈�: �W:�9!�޹r��K���y[�P���������Ň�s����U�K�(��g��ɇ����~��x   x   1�����_�T9����@�޹�f�9=2H:�b�:S�:Vc�:3H:�e�9Ҙ޹��`9���_�:���J\û����
��\���)�K�2��x5�I�2���)��\���
����N\ûx   x   �P����_�������Y߹��c9!,:OWf:Wf:),:a�c9BV߹���x����_�}P��Z�ǻ�7�����*8&�?<7��nC���I���I��nC�B<7�18&�����7��a�ǻx   x   ����&}[�������� Z��+9�:� :X�:�/9�X乧������|[�����K�ǻ:��y6�]z,���@�x�P���Z��!^���Z�}�P���@�fz,��6�-��?�ǻx   x   �����S��	��w��3�����7�ݎ9���9���7����w����	��S�����_û�9��;7���.���E���X��f���m���m��f���X���E���.�<7�:��"_ûx   x   �����|G��S�n������4��>z(���<������|S��|G������	��S����+|,��E���[��m�cx�d�{�nx��m���[��E�<|,���%��
��x   x   ���G�9�������a��a[���\��ێ�Ӛ��ރ��l�9�����e��8�້�
��;&���@�Q�X�-m���{���������	�{�Bm�H�X���@��;&���
��໴e��x   x   vp� �*��M庳����&A�D(��%A�t���#N�;�*��up�U��Kл=���a�&A7��P��f�Ix�e����r��d���/x��f��P� A7��a�N��RлU��x   x   Y�]����غ]���ol��pl��\��%�غF��Y�+ґ�ʠ��eO�J����)�uC���Z�wn���{�-���2��� �{�vn���Z�uC��)�,��RO�格��ё�x   x   �B�JH�'GϺ�ן��֏��ן��GϺ�H���B��Ӂ�O�}!ӻ�!�[���2���I�{)^� n�zx���{�Ux� n��)^���I��2�j��"�g!ӻ`��Ӂ�x   x   1H-��`�f�ɺ�ث��ث�,�ɺM`��G-��Yd��$�����1㻶��!���5�H�I���Z�}�f�!"m�G"m���f���Z�E�I���5��!��� 1�����$��<Yd�x   x   ��*:�Ⱥ>��0Ⱥ�:����G��Q~�~w����û׏��}
��"���2� yC���P�nY���[�QY���P�yC�c�2��"��}
����ûhw���Q~�G�x   x   b	���eUɺEUɺ�⺾a	�}�,��jY��\��W⥻ҡǻ��뻸������)�_G7�x�@��E��E���@�WG7���)��������뻠�ǻG⥻�\���jY�G�,�x   x   �J��A1׺*W̺2׺�K��B��܌8�7�b�(+���㥻�û6��%�d��9h��C&�w�,�ڪ.���,��C&�!h�S���%�+6�.�û�㥻I+����b�Ɍ8����x   x   I�ẹ�ϺӶϺ#�����C�٪<� c�]_��U{������)ӻ
Z���e�
���qA�iA�����
����Y컏)ӻ���[{��6_����b�/�<��C����x   x   u"Һ,�ʺ$Һx��,�E�?�8�lpY��Z~�+��l���i���л������VM��'��qM�����X��5лj�������9+���Z~��pY��8��D�<���x   x   PoȺnȺ �Һ��级��p����,�hG�fd�܁�ܑ�Va���s����qû��ǻ��ǻ)qûM���s��1a��	ܑ��ہ��ed�[G���,��������)�Һx   x   ����٦�&��s����)���?��۴ͺBXܺ���s���	p�"������7�,��Q� �*��J7������hp�K����캀Xܺ��ͺ	?��;*�������&���٦�x   x   �ئ�/����襺�����J���^���>��f����B������}#ʺ�@Һ�-ٺ�?޺��}�ຢ@޺�-ٺ�@Һ�#ʺ����A������l?���^��rJ��[���-饺���Yئ�x   x   �"���楺:���k��?������bӅ�6悺4䁺�x��]���텺8����ڈ�QN��&و������%��{x��L偺�悺'҅�
������yk��꩟��楺X$�����x   x   c�������h��8���r���T��?:��Y$�i��F�����Mz���c��_�f�gg��w��͛�����{��=W$��?:���T���r�Z7��h�����܁��W۴��ܴ�x   x    ��B�������r�b^B����~�ҹ����.�Ս���簶�'8�rz8���8S�z8� 8�=��?����-�;��=�ҹ����\B�}�r�����A��/ ��Iº[�ź�ºx   x   �1���Q��̤���T�{����������*�8k9��9��9���9��:R�:Ӈ�9*�9��9�k94)�8���`�������T������Q��U1��yӺ�rܺKrܺ�Ӻx   x   P�ͺr-��#ą�[':��sҹ�}�f�9�_�9�:@64:��L:�Z:CZ_:��Z:��L:�64:b�:C^�9Τ9Hw�-vҹD':��Å�!-��Ģͺ��j����~��]���*��x   x   %Aܺz屺�҂��8$�j뉹.��8p�9n�#:��W:�~:�s�:
|�:�}�:�t�:�~:F�W:A�#:�p�9��8�뉹7$��҂�o決:Aܺ9���?��5������j���x   x   |�o(���́��c�����|k9��:��W:.i�:�ƚ:?,�:��:n*�:�ƚ:j�:��W:F�:k9���#d��́��'�� {�4=����'��X+���'����<�x   x   ͒��)s���]�����oQ��[C�9hL4:�'~:+ʚ:]#�:ZQ�:�Q�:�$�:#ʚ:&~:!M4:!C�9�V�����\��tr������7����/�?��*G��*G��?���/�,��x   x   [^�Yʺ6탺�2�������[�9��L:O}�:2�:�S�:dȻ:�S�:�0�:�}�:D�L:k[�9�o���1���샺ʺ�^�Y)'��~B���W��d��_i���d���W��~B�h)'�x   x   �v�Һ�ͅ�u���.8���9!�Z:n��:s�:NV�:�U�:��:���:��Z:��9r58����ͅ�7Һ�v��24�[&U��/p�[���>�������l����.p�&U�f34�x   x   %��/ٺK���B��}8�!:�{_:7��:H3�:A*�:�3�:䉑: y_:]#:޹}8V��.���ٺ����?�B�f�^ꃻ�ǐ��똻v����똻�ǐ��ꃻ��f�9�?�x   x   t"��޺귈�I��2�8�":��Z:؁�:uК:qК:F��:4�Z:�$:�"�8��빱����޺�"���I��u�\���ڞ�u����������(u���ٞ�"�����u���I�x   x   �����X+������}8h��9��L:m2~:�s�:	3~:�L:��9��}84�빪*����ປ����P�����Z��A��nJ���û�Fǻ�û�J�����pZ��饀���P�x   x   '� ���Ƕ����\8;j�9Y4:h�W:��W:VY4:}i�9tj8���$���E���� �?_T��Z�����cz���[ǻ��Ի��ۻ��ۻ��Ի�[ǻZz������Z��@_T�x   x   Ȯ��޺ہ��P��dE��FX�9��:��#:�:�W�9Zݗ�S������d޺���`T�����l堻�x��T�л���z�컝��������л�x���堻�����_T�x   x   $��
ٺ[υ��-��U��\�k9ԙ�9���9�k9U��T-���΅��
ٺ�$��P��[��"栻o���5�ջ�Q껳+���v ��v �^+��3R�X�ջ���栻�[���P�x   x   ��u Һ������=�8�9	2�8�|�����탺� Һ���U�I�0���)���Cz��C�ջN.�݌����y��H������.�`�ջ�z��顝�姀��I�x   x   z��ʺ^���^��щ�-�渾���щ��^��]��ʺz��@�Тu��]���}��g�лST�=����b��[��[��b�m���]T�4�л�}��^����u�T@�x   x   zb�Mv���́�/$�3Wҹ�n���Vҹ�/$��́�qv��Ab�j84�^�f���������`ǻ�⻴/������\��U��\�����/�����`ǻ�������N�f��84�x   x   b���l+���҂�5:�W�����:�G҂��+��^���6/'�>.U�B�ߞ��P��2�Ի��커y �Р�o]��]�۠��y ����J�Ի�P��iߞ�fr.U��.'�x   x   ��>鱺������T�HIB���T�o��鱺���+��ņB�:p��͐�@|����û��ۻ���Tz �t��*e�7��gz �����ۻ��û�|��+ΐ��9p��B�h��x   x   eHܺv0��;���S�r�?�r������/��9Hܺ�B��/�D�W�麁���L���Pǻ&�ۻC��64������ݔ���4������ۻtPǻ5���C�亁���W��/�~B�x   x   .�ͺ�S�����$1��d��JS���ͺ����!�c&?���d����q�������� Ļ_�Ի��:\�
7��[껞⻬�Իr Ļ}�������-���,�d��%?�"�����x   x   )6���B���e��Re���B��s6�����y��ֿ'��6G��ni�a����������V���gǻ��л/�ջ)�ջ��л�gǻV��E�������<���zni�7G��'�@�����x   x   {$������G���d���6$���$Ӻ8�� �	d+��8G�i�d�����Ґ�7垻�����������F���؄��|���l��W垻�Ґ�������d��8G��c+������%Ӻx   x   p���祺y楺Ƅ���º�}ܺ���� �C�'�;+?�ܡW�Cp��������f��U�����]�(���g��8�������UCp�ѡW��*?��'�!�W����|ܺ�ºx   x   \%��Y���B&��<ഺ��źܺ�����k'�ş/�W�B��:U�N�f�G�u������f��0����f��᱀�`�u���f�!;U�$�B�ǟ/��'�������~ܺl�źഺx   x   �٦�W٦�&����ⴺMº�*Ӻ��纏���J�_���;'��G4��@�g�I���P�vT��uT���P���I�A@�KG4�8;'�����J��
��o��?+Ӻ�º�ᴺ[���x   x   N'��
������T��?i��|釺����Q�����ᇺ�>������&��hq��m����͉������p��P��T����>��Eㇺ����K���`���_臺{j�����>���
��x   x   �	��"D������������v�ݴk��`�hV��hL� �C��=<�)6�CZ1�W&.��y,�|z,�@'.��X1�T6�2@<� �C��fL�tV�ܟ`��k� �v����������C��
��x   x   �������L�{���i��U�W�?��%*�_��ۀ�W����ʹvt��������­��E��!��1w��w�ʹ����x���!*�Ԁ?��U�|�i���{�����웉��>��x   x   �������̍i�%HM��8.��T�c�޹�ݤ�۾b���	�xQ��%C���:�7RJ8�/J8�,�7�[���V���
��b�Fڤ���޹AY�~8.�GM�G�i����#��Ip���p��x   x   �d��C�v�
U�&5.�U������BN�t]v�P��8��*9�~9�Q�9�-�9���9�/�9�P�9C�~9"�*9���8�Uv��HN��}��5��+6.��
U��v��d��1����g�����x   x   �⇺=�k�kw?�rL��w���/$�x��7��?9�է9��9�6:�D:��:b�:rD:�5:��9�ק98�?9/��7�-$�Py���N��v?��k��⇺ݝ��G-���,��c���x   x   ҍ��э`�,*��޹FN��(�7Dk9Q�9�:�#.:d�C:�%Q:{�U:�#Q:<�C:z$.:;�:�P�9�Ik9�M�7#N��޹�*��`�͍���O��+l��q5���l���N��x   x   w��t�U�?������K�u�u@9!Z�9�H:�/B:L?`:�Gt:G~:�H~:�Gt:�=`:�0B:�I:\Z�9>@9D�u��������U�zw�����ɼ��b"���!������+���x   x   r����NL�{h��hb�"J�8��9��:;4B:�i:��:��:d�:v��:��:��i:	4B:��:��9�]�8olb��j��ML������������HǺ �˺*HǺΪ������x   x   c҇�ʟC��N湷�	�
+9�;�9�0.:MG`:��:Yʏ:��:��:�ʏ:��:�E`: 1.:w<�9�+9F�	�sL�ޝC��Ӈ�Gw����ĺ�غB����ẜغ��ĺ�v��x   x   K-��<�ԋʹ�n���V9K:D:�Rt:��:q�:���:_�:���:RSt: D:�J:TW9j����ʹ�<�P-���Ǯ��Ϻ������i�������W��(�Ϻ�Ǯ�x   x   q���9�5��/����鶷��9)[:�7Q:�T~:�h�:��:��:zi�:�U~:S7Q:�Y:"��9ۏ� 1����5�H���R����ٺU������J��K�&�����ٺ`���x   x   y����21��գ��_�7�g�9U	:��U:�X~:A��:�Ώ:盋:�W~:��U:�
:�k�9/M�7�գ��21�����k��d[��4��t�q���`p�`u�I6��Z���x   x   �[��X�-�]ę�G~L8�ط9�:�9Q:QYt:Y!�:�!�:|Yt:�:Q::kԷ9?qL8ę���-�}\��s���)b뺚�Yv��(�	N/�EN/�!�(�bu����c뺩���x   x   7����O,�m_���jL8�n�9�_:�	D:�O`:��i:P`:9	D:R^:�p�9�L8]���P,�˝���2�����*���%�U�4��>�BSB�=�>���4�N%�I�����S2��x   x   I���:P,�k�����7���9\Q:�;.:OCB:dBB:�;.:mR:��9���7�����P,�~���∿�׀����J�+�j�>��[L��nS��nS��ZL�e�>��+����������x   x   ����y�-��ң����t9GR�9�:\:��:>Q�9�t9�7綱У���-�����9��������	�/���E���V���a�	9e�q�a�:�V�{�E���/�2����������x   x   �[��T01�K+��fA��y@+9��9�|�95}�9��9�<+9_7���)���11��\���3���������a1��I��e]�B�k��
s��	s�y�k�f]��I�a1��������J3��x   x   �����5�~ʹr	�k��8V@9D�k9�Q@9���8߀	�;�ʹ��5����������R��M�/���I���_���p�E�{�,��Q�{���p�ͭ_�ĀI���/���������x   x   ����4<��B湑Cb�*�t�)f�7ߒ�7w�t��Fb�=A湲<�ϗ��v���e�W����+�W�E��g]���p�7�~����I����~���p��g]�*�E�D�+���f� ��x   x   �-��R�C�;d�M����M�Y�#���M�����d�G�C��-�������_�l�%�+�>���V���k���{�F��Є�M��\�{�]�k��V�l�>�[%���_�G���x   x   ;ԇ��IL�	���k޹T��oX��:l޹{���JL�^ԇ�4ʮ���ٺE8��z�2�4��`L�Ύa��s�Q����������$s�<�a��`L���4�)z��8��ٺ�ɮ�x   x   ����)�U�}
*��D�T��B��*���U�&���z��تϺ�$���y���(�k�>��uS��?e�Qs��{�p�~���{��s� @e�QuS�`�>��(�z�C#��{�Ϻ�z��x   x   �w����`��m?�(.��).��n?�1�`��w��M����ĺF�躦��3w�'U/�([B��vS�ڒa���k���p���p�
�k�X�a��vS��[B��T/��v��������ĺ����x   x   䍇��k��U�';M�IU��k����ƃ��+���غ���#Q�#���V/���>��dL���V�fo]�O�_�1o]�v�V�HeL�A�>�=V/���QQ�G���غ����Y���x   x   �ᇺԲv���i���i�"�v��⇺TR������lOǺ��	���R�y���(��4�%�>�5�E�*�I�@�I���E�l�>���4��(�y��R��	����
PǺ����R��x   x   f��ڈ���{�R����d��
����p��])����˺�
��������~����%���+�-�/�l1��/�R�+� %�����~�H�������
��˺)���p������x   x   ����������������,1���;���*��ZSǺ?غp�躐-���@����f������b��c��J�~?��.��E��1غ�SǺ�*��w<��f0��Ξ��x   x   �����B��қ���q��k���1��nt���Ʈ�P�����ĺ]�Ϻ]ں�o�kz�4��������F������Fy뺨p��ں��Ϻ��ĺ���7Ʈ��s���1���l���q��x   x   �	�� 
��W?��&s���������?W��
�����5����ٮ��Ƴ�>"�����jI��c���럿�bI��񶻺N"��{Ƴ��خ�M����������X����������r��n?��x   x   %�a�t$`�}�[���T�v�J�Α>�e�/�oO�ޫ�!G��r0Թ賹�N��3���k�V�b�e�k��3���P��賹w-Թ�J�����LO���/��>���J��T���[�s$`�x   x   �$`�"�[�]nS�VG��(7��i$���Ѣ��^Ź���#`��J�����W�8��ɻ�.�W��༸�I��*`�E���\Ź���v��l$��)7�G��mS���[�h%`�x   x   ]�[��mS���E��3��������Gҹ�����M�2ѸQws��m8L�8s�9M�"9z�9�>�8��m8is�+zѸqM������Dҹ���y��V3��E��mS���[���^�x   x   ��T�	G��3����������t�z�e�����춮P�8��@9�9�V�9M�9N�9�X�9��9��@9�H�8�"����R�z�#���������43�G�0�T�j�[���[�x   x   �J�@&7����ӽ��n��0JZ� ᔸ�F{8y�<9Ý�9��9�(�9�5�9� :�2�9�&�9��9ԝ�9��<9)X{8�甸$GZ��i��9���D��	(7���J��,W��H[��-W�x   x   ō>��e$���>�BZ��?b���8��u9�i�9%�9��:Bq:%:%:�r:!�:��9�j�9Y~u9��88Bb��FZ�6�d��>f$��>���P���Y���Y�;�P�x   x   ��/����;ҹ��z�Y�%,�8���9f4�9a�:j	":E�5:r�A:��E:5�A:��5:
":I�:r5�9���9�0�8`���=�z�S9ҹ����/��5H��aW��\�%bW�3H�x   x   �G�a��Л��h��O�{8>�u9�8�9[�:�,:�cD:eU:i�]:̪]:�U:�cD:�,:��:�8�9�u9G�{8�b���ћ�\��KH�[�=��AS�^B^��B^��BS��=�x   x   ��vJŹ��L�4O�H�<9>v�9��:�,:�kI:�_:�^l:�p:N^l:S_:	kI:!,:��:Uw�9�<9ב���L�lIŹ-����1���M��^��d�ջ^�,�M��1�x   x   �/��_��) Ѹ���8���9�"�9�":&hD:�_:)Vq:��z:�z:�Uq:_:8hD:�":�#�9���9��8jѸ���3��i�$�3CF���]��i��i�i�]�5BF�/�$�x   x   �Թ��_��p�ܸ@9H3�9ڑ:��5:� U:�bl:��z:�]:x�z:�bl:� U:6�5:Ñ:T4�9.�@9��o�5�_��Թ�r��=�E�Z�,m�#Bs�um�7�Z���=��r�x   x   'ɳ�Z�B�n8��9D�99}:��A:��]:!�p:	�z:f�z:��p:�]:P�A:�}:_B�9_�9��n8	��ȳ��C
���4���V�x�n�LV{��W{�S�n�
�V�߶4��D
�x   x   M,���a����8�w�9FT�9�!%:��E:��]:fl:C[q:�fl:ų]:Q�E:�!%:(U�9�w�9<��8d��\*��������+�p/R�R[o�mЀ��胺�π�f[o��3R���+�����x   x   ���lyV�.�9q�9� :R$%:��A:D&U:�_:W_:!&U:��A:#%:ʹ :!r�9?�9HrV�#������#�3aM�g�n�XL��n��9n���L��3�n�^M���#����x   x   �mk��o�K�"9�t�9�V�9|�:��5:dpD:�uI:�pD:��5:C�:�Z�9�t�95�"9�p��jk��ڹ�z�:I��Hn�\V��@��}E��0@���V��Kn��I��x�$�ڹx   x   �Sb�#h���9���9<M�9��:�":o$,:�$,:D":&�:�M�9o�9��9�_��Wb�Bhӹ�t�VF�e�m��݆�t0�����p��g/���݆�2�m��F��w�iӹx   x   ek��CV����8��9�C�9 7�9��:��:��:�7�9wD�9��9_��8BV�dk��fӹ��t�D��'m�出�,��m���n��鐝��-���䇺D*m�P�D���hӹx   x   ���T.���Ko8��@9�ŕ9���9CV�9LU�9���9�9��@9�So8�=������ڹ�s�=�D���l��g��e���~���禺�妺�}������g����l��D��u�Q�ڹx   x   :%�����c�m����8Q=9�u9۲�9��u9�$=9���8G�m����!����蹸x��F�
(m�h�����0���8��ܕ��T
��l���N����g��)m�F�Gv�r��x   x   ����e�_���и���܋|8m��8���8Mm|8���*�и.�_�g�������_�#�?I���m��出�������s���������r��,�������出�m�I�k�#�����x   x   9Թc򘹫�L�\	��LW���=a�QM��4����L�8�Թ_?
���+�`M�eIn��ކ�.��i����	������4�����i�����~-��R߆�-Jn��]M�A�+��@
�x   x   �%��97Ź�����z�BZ�8Z���z�e��� 8Ź�%���m�ε4�E.R���n�}W��B2������
ꦺ8������������馺璝�2���V��U�n�/R�3�4�lm�x   x   ��҅�#ҹrڼ��L��׼�
$ҹ���w����$�=�=���V�-\o��M��TB������q���馺����u�����Gꦺ�q������B���M���\o��V���=���$�x   x   A��v����¥��2���"���w��A�k�1��@F���Z���n�
Ҁ��p��I�������������8���w���M���_���<���I��"p��]р���n�,�Z�@F�+�1�x   x   �/��_$�����׼��^$���/�r�=���M���]�m�"Z{��냺1r��	E���4���3�����U���%��?2���5��qE��sq��6탺�Y{��m��]��M���=�x   x   ��>�0 7�C3�3�M!7��>��2H�d@S���^���i��Fs��]{��Ӏ��Q��]��E䆺�뇺�n��o��P쇺C冺�[���Q���Ӏ�N\{��Hs�ʥi�ֿ^��>S�2H�x   x   �J�7�F�|�E���F���J��P��`W��C^�6�d��i��m�Yo�]fo��n��Yn���m��:m�`m��9m�u�m�WXn���n��fo��o��m�P�i�d�d�5D^�*bW���P�x   x   ��T��iS��iS� �T��*W�]�Y���\�JF^�H�^�դ]���Z�v�V��@R�mM�<,I�S#F���D���D�S$F�v,I��mM�z=R�g�V�%�Z�y�]���^�wF^���\�3�Y��)W�x   x   �[�[�[���[�'�[��H[�3�Y��eW�CHS���M��KF�U�=�;�4���+�i�#�������V$�ȉ� ����#�0�+�|�4���=��KF�@�M�vES�]fW��Y��J[���[�x   x   �#`�U$`��^���[�./W�Q�P��7H���=��1��$����S
�y�����L�ڹ(�ӹ��ӹ{�ڹt鹑����S
��_�$���1�f�=�B:H�Q�P�-W�9�[��^�x   x   I�2�b�0�*�+��["�Y����O�ݹ���F�t��Q
�,�v�y8F�9!P9Z�w9���9.�w9)P9��9��y8n�eS
���t�H��S�ݹ`�� ��\"��+�^�0�x   x   ��0�7�,�4&$���5����๖��|Qu����՞��"��8b�,9a�w9��9��9ό�9r�9��w9N�,9���8Ѻ�q��7Vu������๝�����%$�P�,���0�x   x   �+��&$������j;��2���r�Hk��J,�6��8��J9Z�9>��9��9ם�9;��9���9��9%�J9���8���e���r��3��j6�ۓ�����&$���+�.�x   x   �\"�G �����e⹔̯��on����~�_6�/�8��g9���9���9��9#o�9�s�9G��9��9��9�g9[*�8 �]6���on��̯��i�X����3]"�)(��(�x   x   P����d;�O̯�_�l�㸎�R7e
99�9Io�9cg�9_� :!:�:+:@� :se�9p�9o�9
9{S7��z�l��̯��6⹊��,��m�#�!�ao�x   x   ���3��P2��-nn�N�Vn�79�ԇ95��9���98�:�C:�=!:�=!:YF:>�:L��9���9�ч9�9�c�7&�mn�3���๹����?�����n
�x   x   s�ݹ:���r���츞1S7M9��9Rb�9]>�9Y:��%:cu0:4:�t0:��%:�:�=�9�c�9s��9�9�S7����r����%�ݹM���ɏ
��&�%�
�����x   x   ��Ou��a��Za6�
94ׇ9�c�9�� :�s:�L-:�(;:BRB:�RB:k*;:M-:|s:m� :�b�9�և9�
9�[`6�e���Lu����׹ƅ��
����׹x   x   Y�t�������A�8��9}��9�A�9�t:�/:��@:�JK:}�N:�HK:u�@:Z�/:du:�A�9���9Z�9�@�8�t����+�t�����{˹��q�&��}˹����x   x   �N
�nd��P��8��g9�u�9���9$:�N-:��@:�kN:��U:ӏU: kN:f�@:�O-::��9�s�9��g9���8t���N
�R�m����� ��gDȹ�KȹA"������`�m�x   x   ��uʡ8K9c��9]p�9��:��%:<,;:PMK:�U:7Y:�U:NK:?,;:�%:<�:�p�9���9�K9'ġ8-��D��k]�ӎ�g����[�������Ԏ�o]��B�x   x   �z8��,9�(�9���9*� :�I:�z0:-WB:��N:��U:��U:��N:�VB:xz0:FK:� :��9�%�9�,9Gz8���K��b�B�C�r�����*����r��B������ �x   x   ��97�w9���9u��9J:�D!:4:&YB:TNK:}oN:QK:FXB:\4:?D!::���9��9z�w9I�9XE8�z�}�Ѹ����.=��3H�O.=�I��РѸ_���lE8x   x   "%P9��9>��9I�9��:,F!:B}0:>2;:Z�@:�@:�0;:[}0:�E!:+�:с�9 ��9D�9$P9$��8qI.8.����>����޸���E��
�޸'>��^!��p>.81��8x   x   <�w9���9���9���9*:jP:N�%:8V-:��/:�V-:��%:~O:�:���9���9@��9��w9��,9(�8�58�'N����s�J���s����\YO�� 58-9�8�,9x   x   �΂9%��9��9ح�9�� :|�:g:�}:�~:�:�:[� :1��9z��9���9�͂9gG9"P9!ֻ8�pT8���7�+�5<��+����56��7�T8Gڻ8�G9hG9x   x   ��w9c"�9㚰9
��9~�9��9KU�9�� :�U�9��9[��94��9���9? �9��w9glG9�t9���8�S�8�τ8�^H8�- 8�8� 8rHH8̄8�P�8���8`{9�hG9x   x   �2P9(�w9T4�9���9n��9���9}�9[z�9E��9G��9���9�4�9�w9�8P9�,9`Z9���8�9�8F%�8�*�84��8�v�8���8��8�0�8�%�8�:�8���8�U9]�,9x   x   95-9�+K9$�g9�9x�9QƊ9X�9��9��g9.K9p-9e9)�8|O�8^�8�f�8=.�8�g�8�`�8��8�k�8ƚ�8�Y�8�e�8h1�8�a�8s��8�\�8��8x   x   ћz8r�8�E�8���8�U
9	Q9�O9N
9��8y=�8��8�z8��E8M�.8p{58�T8�8�:�8�g�8q��8�[�8�b�8��8al�8�5�8��8u�T8�i58��.81�E8x   x   KZ��>��3��M`k6�zV7��7%�V7��l6@����)k�'m����������G�k,�7��H8$8��8�_�8���8�]�8���8dɖ8��H8�	�7&H��D�����T|�x   x   x&
��������Z�2��i��<^�3��s���$
�X�!���\JѸ����#�ҥ5�m 8t��8x�8h�8_�8a��8��8�Z 8`��5��I���VѸ����"�x   x   +�t�;(u���q��>n��l��=n���q�]!u���t���m�F]�.�B�L���޸J@s����!Q8w��8���8
�8���8 ��8>8����\s�o�޸N����B�G]� �m�x   x   !������������������� ��n��֪��}��������r��=���������3I 8_ʖ8"_�8�j�8�Ö8�L 8����������=�F�r�TĎ�[z��:���x   x   ܜݹ0���#��V�K$���์�ݹ��ֹ�j˹$��>���S����H����Xs�a��51kH8�7�8�c�8	-�8уH8��5/vs����H�~��ƨ��7��0k˹��ֹx   x   ���L��/�����޺�:�������w�A�27ȹO��s����=�U�޸�]���7ӄ8"�8^%�8uل8=��7>D�X�޸�=������S���9ȹw��s����x   x   ��������3���
�l�Xf蹜Aȹ^�����r���H)����M�E�T8]J�8m*�8AH�8��T8�L�*7��r����r�W����<ȹ+b蹼�C�
���x   x   YY"��!$�<"$��X"�Ni�����"��q�1���Ύ��B�@�Ѹh����48pλ8y��87��8C˻8
58i����Ѹ��B�Oώ������<� ���Bi�x   x   ��+�ؾ,�#�+�.(�#�!����V�
����!y˹����i]�H���
��/.8C(�8Y:9�h9�=9g$�85.86u�N ���f]�p����v˹�|�0�
�t���!��(�x   x   ��0�q�0��.�(��m���s���x׹����C�m��B����PE8ػ�81�,9!SG9fNG9�,9���8�UE8D��A���m�!���N׹�����k��(�".�x   x   �e�s���%�7\��ӹ����77���J �o�C�S��8�49�Ҏ9�9���9�A�9`��9wC�9`|�9��9�ю9p�49���8��C�VI �s7�������ӹ�]�%�i��x   x   ��5���)��Нܹ�c���!��?�C��
�����7W4	9�nt9���9�d�9^��9m��9��9���9yf�9sĩ9mt9.	9��7'��b�C�.#���e��_�ܹ)��ˠ����x   x   �&��*��O߹����?=��:�X��下��5S�8m�W9Nt�9hq�9�w�9^��9.:(��9|x�9�l�98s�9��W9~T�8:�����N�X��:��o���uS߹_*���&��Z�x   x   �_��ܹ����ො�L�b������ڨ�5˲8Y-F9b��9���9!��9A :�:
�:� :���9l��9���9�,F9>��8TӨ�d����b�.���������ܹ	`�P�������x   x   ��ӹ�f��1?���b��$�$巢Ο8+�<9�4�92#�9���9>G:�:"�:2�:�F:>��9�#�9�4�9u�<9�џ8�#�$$�E�b��<��|i��L�ӹ��⹵��@��x   x   ����,&����X�������&�8��89ӫ�9�E�9���9!�:ѩ:��:��:׫:@�:֖�9�G�9騐9l�89o*�8O州���[�X��'������k�ù�ι�ιB�ùx   x   T>����C��)������ʟ8�89K�9v��9�I�9��	:+�:�� :��#:�� :.�:<�	:G�9{��9�M�9͋89z̟8�����*�ٛC��>������J���r��%K����x   x   <[ ��"�� 	��w��8�<9���9���9T�97�:.�:;�&:ݵ,:��,:��&:S�:6�:`U�9a��9𢡄9f�<9潲8e��!���Y ��X����\���߼��>����X�x   x   ��C�$Z�7:B�8�(F94�9)F�9�J�9��:�:OQ*:˲2:M�5:A�2:SR*:L:�:�J�9DF�9�4�9�'F9�E�8�\�7	�C���ٸ�]�>�4��(>�(�4��_���ٸx   x   H[�8�&	9U�W9���9i#�9��9��	:R�:R*:��4:�.::%1::a�4:�Q*:K�:��	:D��9�!�9���9�W98%	9�^�8��6�}�a��@���0���g���m�b��6x   x   %n49:bt9�p�9��9@��9��:/�:R�&:��2:�/::��<:�/::��2:�&:?�:�:��9"��9�p�9�_t9�n49T:�8Dc�8��<8��7�&�7�k�7�<81`�8b@�8x   x   �Ɏ9&��9co�9��9�H:b�:�� :�,:,�5:C3::�0::<�5::�,:%� :ѭ:�I:h��9�k�9���9<ˎ9��n9@�G9��)9��9jJ9=H98�9��)9�G9�n9x   x   >ۻ9�`�9^w�9� :��:c�:��#:�,:L�2:��4:�2:l�,:�#:m�:�:� :�w�9}c�9�ػ9j$�9q��98i�9�g�9ࠃ9�9%��9Zj�9�f�9���9w&�9x   x   �{�9j��9M��9��:)�:��:9� :��&:�W*:�V*:��&:�� :��:��:j�:ֈ�9��9�y�9(��9���965�9!a�9&+�9�"�9�#�9<*�9_�9(9�9���9+��9x   x   ,>�9��9U0:�:��:�:��:�:�:��:�:��:��:��:0:���9?�9�z�9}�9�|�9.��9hL�90�9}��9@/�9�M�9���9qy�9�#�9�y�9x   x   ���9}��9���9� :@M:��:%�	:�:x�:��	:��:�N:z :P��9���9ݹ�9Kh :qT:�	:��:��:n�:��:��:��:��:_�:G	:�S:�h :x   x   �E�9$��9҂�9G��9���9��9�X�9!g�9y[�9��9A��9���9���9���9�D�9�i :3V:�F:n:(�":T�):.:Π/:�.:�):��":�n:+F:W:�i :x   x   Ӂ�9�o�9�y�96��9�5�9�Z�9��9���9�X�9e3�9���9�z�9�p�9��9���9�W:�H:ʱ:6r+:k36:+�=:�B:^B:Z�=:Z46:Lq+:m�:HI:"V:���9x   x   ��9�Щ9~��9��9QH�9z��9�b�9���9�H�9{�9b��9<ϩ9��9���9�*�9�	:eq:�s+:k|::~5F:��M:\3P:��M:�4F:}::�s+::p:	:,-�9~��9x   x   �܎9V�t9�X96SF9��<9L�89U�89ȸ<9�RF9X9��t9�ގ97�9��9���9 :5�":�66:*7F:ťQ:��W:
�W:�Q:�6F:�66:k�":B :���9���97�9x   x   ��49=M	9���8��8_&�8���8�$�8!�8ޞ�8�Q	9)�49
�n9h��9�H�92��9��:׵):��=:�M:�W:�[:�W:��M:_�=:״):�:���93M�9M��9�n9x   x   $��8��7�������n��o�㷙���݀��R��7��8���8��G9��9�v�9�`�9��:�.:�B:�7P:��W:�W:b7P:�B: .:�:c�9�s�9�{�9��G9��8x   x   v5C��Ұ�.��kv�����Wz��)�㸢Ȱ�W@C�{��6Aà8~*9��9fB�9�E�9o�:H�/:'B:��M:y�Q:��M:WB:��/:��:�B�9�B�9X��9�*9�Ġ8�J�6x   x   �. ��oC���X�0ub��ub�%�X��rC�/ �5jٸ����=8K�9g��9�:�9��9��:� .:~�=:	:F:�:F:��=:,!.:Q�:���95<�9���9"�9И=8����eٸx   x   z+��|���+��'����+������+����X��2����Z��7{9G�9J;�9�E�9��:��):\;6:M�::n:6:��):�:"C�9�;�9c�9�}9~��7f��^5�}�X�x   x   놯�Z������ڽ���Z��焯�����a�Х4��ï����7�v9D��9�@�9�b�9��:��":�w+:Ix+:Y�":Y�:�c�9B�9H��9�{9WS�7�̯�!�4��z�����x   x   ��ӹ�ܹ�H߹!�ܹ��ӹk�ùz;��b����>�᯸���7��9��9�s�9D��9�:�u:��:�s::i��9ir�9���9��9��7�ӯ���=�����}>����ùx   x   SX�"��V"���V�"��ι�e������T�4�!���t=8��)9}y�9�J�9��9�	:BK:�L:�	:��9�J�9{w�93*9l=8�����4�����#a���ι9��x   x   T#�q���#�V���n��-ι�?��Ő�bC�2��R��8��G9ֱ�9���9�/�9>X:?Z:�W:�,�9���9���9,�G9���8���JD�҆��B���ι��繯���x   x   ���9���X�����ؿ��ù����ԺX�o�ٸ ��6(s�8էn92�9B��9y��9gk :�j :n��9$��9m0�9s�n9�q�8}��6Ԑٸ!�X������ù8�⹔���0Y�x   x   �+ƹ`�¹,��x5���a���0U�k)����I�8��59[�9�K�9"|�9��:�@:��:x@:(�:>|�9�K�9��9��59�F�8��3-�70U�/c��i6���*��B�¹x   x   ��¹PV��-����M���p��&�0���~�7D��8Qb9	ۢ9'-�9�B�9`:�:w�:Qa:�D�9r.�9bآ9�Ob9Y��8~X�7g/���&���p�3L������X��n�¹x   x   �.��b����o��f�}��y:��Ըނ�*ˡ8˩49c��9R��9���9���9J�:p�	:�:���9���9���9A��9��49M͡8 ʂ���Ը_|:��}��q��⠬�<-�����x   x   V9��PP����}�R�@��(�4���+a8�z9v9B��9���9פ�9��:;Q:?R:��:��9���9���9�v9�{9�-a8¬�g&���@��}�nO���9���<��M;��x   x   �f����p��~:�:-���#���48j�9�uc9�Ý99��9R��9�� :g�:�:c�:%� :��9���9QÝ9yc9��9�48��#�l/�Ɓ:��p�h�����P���G���x   x   �>U���&��ո[��Q�488,9�x[9���9�M�9_��92� :��
:��:��:��
:�� :��9�P�9���9�v[9C19��48����ո��&��<U��t�����P�����t�x   x   a;�7L��0���a8��9Uw[9�9���9���9�<:��:&:(�:�:�:�=:���9̮�9	��9iu[98�9a8u+���L���=���'�F�>��[F���>�ح'�x   x   ����7��8�r9$qc9���9���9/��9�:Z�:r�:c:�b:��:�:��:���9B��9��9�sc9�u9���87ߒ7���n&��]�̸[��݊�:�̸r,��x   x   �8��8��49��u9���9�L�9���95�:8s:��:/\ :W�":�[ :h�:>r:&�:$��9�M�9���9@�u9�49'��8�8�Q�7���5d������vW����5]e�7x   x   ��59�;b9���9l��9���9��9�<:��:'�:��!:��%:m�%:W�!:��:��:�<:ɥ�9M��9H��9J�9=b9��59r�9��8
��8[��8B��8E��8���8��9x   x   ���9Т9���9"��9���9z� :��:Ŀ:\] :�%:2�':��%:X] :]�:��:� :ۨ�98��9���9�΢9���9�b�9Wn9w-^9�T9~�Q9�T9.^90n9�c�9x   x   =�9y"�9���9Z��9˺ : �
:�:.e:]�":�%:y�%:��":
e::r�
:�� :���9V��9�"�9�=�9��98o�9�ڮ9e�9�˪9�ɪ9Z�9@ܮ9Kn�9��9x   x   Rn�9�8�9���9��:�:��:�:f:�^ :��!:*_ : f:~�:��:Z�:"�:O��9f<�9�m�9C�9���9���9}��9B��9M�9���9���9���9���9��9x   x   V�:�[:b�:AQ:4�:��:[:��:a�:�:/�::ȷ:��:]Q:f�:\:f�:)�
:�)::�:0{:�:��:�z:��:�:�(:�
:x   x   �;:!�:��	:sS:C�:��
:��:A�::w:�:��:��
:��:�R:E�	:v�:�;:U:� :G�(:ia0:_6::@::Ǚ;:@::X`6:ha0:j�(:&� ::x   x   �:��:��:.�:=� :?� :�C:��:�:)B:�� :�� :��:�:��:p�:ʢ :%�,:�=9:PE:��N:<>V:�Z:�Z:[=V:��N:YE:
=9:G�,:٢ :x   x   &>:9a:���9���9��9���9k��9���9���9߲�9��9���9���9v`:�>:U� :��0:�A:R:�`:��k:�(s:*�u:�(s:�k:΅`:jR:ܬA:��0:� :x   x   v�:�G�9B��9
��9z��9e_�9=��9꼿97]�9j��9���9��9�H�9��:�:c�,:үA:��V:p�i:��y:���:҂�:n��:��:Ƞy:K�i:*�V:Q�A:��,:C:x   x   �}�9.4�9᫷9ŏ�9�ѝ9	�9���9%
�9ӝ9e��9ԩ�9d3�9}�9J�
:?� :�B9:�R:N�i:�S~:�1�:+H�:��:I�:A1�:U~:��i:R:�C9:$� :y�
:x   x   GP�9��9��9�"v9�c9'�[94�[9��c9�v9C�9��9�P�9�0�9V2:C ):,	E:y�`:e�y:�2�:U��:Qp�:�o�:`��: 2�:>�y:ό`:?	E:��(:1:]0�9x   x   ��9�cb9q�49$�9r9�T9T9^�9�49afb9�9j5�9���9g:k0:�O:��k:M��:J�:5q�:w��:2q�:�J�:M��:`�k:KO:�j0:d:���9B5�9x   x   �59��8�8�a87^58,i58��a8��8y�8��59z�9憳9T��9��:.j6:ZHV:e1s:b��:{
�:9q�:�q�:�	�:H��:2s:�GV:	k6:��:���9Y��9�x�9x   x   Ll�8��7쁷�0�?#��3������$�7;s�8�9lNn9=��9_��9�:|L::BZ: �u:���:OL�:���:�K�:䆅:G�u:�Z:cL::i�:��9���9�Sn9�9x   x   �B�� ��X�Ը8����&�Ը���'J����7��8k`^9,�9y��9�
:˦;:�Z:�3s:���:�4�:�4�:��:4s:�Z:a�;:�
:���9�*�9]Z^9���8Q��7x   x   �Cu&��c:���@�"d:�3w&���f֔�P��5z(�8��T9��9�h�9�
:jM::�IV:�k:�y:|\~:ϩy:%�k:JV:mM:::Li�9��9��T9(�8�F�5�ڔ�x   x   T U���p�K�}�֬}�[�p��U���'�eS̸s��]�8��Q9g�9$��9A�:nm6:�O:x�`:F�i:��i:�`:�	O:m6:?�:���9��9��Q9�X�8{��Q̸D�'�x   x   �\��FD���h��E��%\����t���>��A踔x��T�8��T9)�9���9��:�m0:�E:2R:?�V:JR:�E:Bm0:��:v��9�)�9-�T9�T�8�}��VE�]�>���t�x   x   �1��d�������%1��猘�����?F��G��&���8�[^9��9���9p:y):�F9:H�A:�A:�H9:�):�:���9C��9U^9\�8���K�W:F�c���R���x   x   �'���S���'���5��Ŭ��Ά��@�>�Ph̸�&�5��8Fn9���9#��9�2:�� :j�,:o�0:q�,:K� :t2:q��9ꂳ9�Kn9��8�Y�5c̸��>���������5��x   x   ˭¹��¹����5��d���&�t�#�'������S�7r9/u�9�0�9p1�9>�
:c:� :y� ::��
:�/�9�1�9�s�9d�9�a�7�����'���t�����97�����x   x   �+����Tp��\O��� �?�ȸ��׷Df8s�9�w9s��9�-�90g�9J�:�/:U:�.:��:�f�9�.�9!��9�w9^�9�!f8$#ط��ȸ� �E]O�$Tp�����x   x   K�p�v��<\���4�y����	{���Q7u>�8�];9;��9:?�9���9�^�9Y	:!:!:�Y	:Q`�9���9�<�9M��9a;9X;�8�vQ7��z�������4�r<\�W�v��x   x   Zp�H?\���:�x��R����d���{8g�94g9�"�9:h�9G$�9�0�9�v:�#	:�v:�.�9#�9�i�9�#�9��f9��9d�{8(�d�|�������:�>\�5Yp�|�v�x   x   �dO���4�����[��r ٷb�.8v��8Z�H9�>�9�ͱ9	�9���90� :fn:pn:� :Z �9H�9�̱9�>�9��H9<��8��.8��ط0O������4��dO��\�2�\�x   x   )� �(��������ٷ8��8�g89�K�9��9�L�9���9e�9E�:�:S�:��9���92K�9<�9�K�9kc89��8B8~#ٷ��������'� �-�4�{�;���4�x   x   V�ȸ,5{��2e��.84�8�639u�{9oA�9J^�9�}�9{��9@�:��:d�:��:���9e��9�_�9�@�9-�{90939g�8/�.8S�d�&*{�W�ȸ���U�
�+�
����x   x   Ɇط��P7�{8y��8�c89Ȏ{9�|�9�9.H�9~�9r:�W
:>U:�X
:�r:z�9�D�9��9�}�9ď{9_89��8R}{8{�P7M�ط!5b�'��D������Cb�x   x   �e8,�8�9s�H9�H�9@�9��9R��9��9�A:�v:j8:G7:Eu:�A:<�9��9{�9�=�9J�9��H9�9��8��e8;��7��68����e���Y�6��7x   x   n9�I;9!�f9V9�9��9�\�9�G�9��9ɝ:v�:3�:6�:�:��:k�:��9�C�9`^�9��9�7�9��f9�K;9Mp9���8���8U�8��8�J�8ڵ�8Ç�8x   x   hw9�9q�93ȱ9zI�9y|�9|�9�A:��:�:��:��:�:�:lB:G
�9F~�9�H�9�Ǳ9,�9��9�ew9�/_9-JM9}�A9C�;9�;9��A9`EM9O0_9x   x   ���9�3�9�_�9��9)��9���9�r:Gw:��:&�:�[:>�:��:�v:oq:w��9���9	�9�^�9A2�9���9(��9��9C!�97�9}M�9��9�"�9��9+��9x   x   ��9��9&�9&��9��9��:�X
:�9:��:��:��:]�:*9:EZ
:O�:��9���9��9T��9M�9��9*��9
�9I��9� �9g��9I��9x	�9���9n��9x   x   7X�9�S�9�)�9o~ :�:��:W:x9:J�:�:D�:�9:{V:%�:V�:,~ :&�9pU�9�W�9�N:T:��:U�	:<:x�:�=:[�	:��:b:�N:x   x   V�:;T	:�s:rm:x:G�:H[
:Ox:��:��:y:�[
:�:�:%m:�t:2U	:k�:��:�6:�� :)G&:q*:5�,:�,:�o*:*G&:{� :�6:��:x   x   �):+:$"	:�n: �:��:{v:�E:S�:F:�t:�:1�:-n:�!	:�:�(:�� :pI+:A�5:� ?:j�F:�kK:�M:mK:ƙF:� ?:$�5:�I+:�� :x   x   .P:D:Cv:#� :�9}��9w�9��9e�9C�9���9�9� :w:�:�P:��':�6:l�D:SR:��]:�f:�xj:�xj:f:��]:�SR:ͬD:�6:
�':x   x   +:�X	:0�9�9J��9��9�O�9��9�N�9��9Ҟ�9�9d.�9�X	:W+:�':�9:�{L:�y^:Qn:>�z:P�:���:gP�:�z:Qn:�y^:{L:=�9:��':x   x   ��:R`�9�&�9X�9�T�92k�98�97�9'k�9$U�9Z�9�'�9`�9S�:�� :�6:T}L:ܥb:}�v:��:U�:��:"�:��:V�:��v:'�b:0}L:�6:�� :x   x   �e�93��9�o�9�ձ9o��9PM�97��9�K�9��9ֱ9.m�9���9�e�9'�:$O+:�D:}^:G�v:^�:�_�:]��:�i�:(��:�_�:7�:��v:b|^:�D:O+:�:x   x   {0�9�A�9�+�91I�9SX�9ܬ{9�{9KY�9�G�9y-�9�B�9(0�9!W:�>:��5:zYR:BVn:~�:�`�:�ە:UÙ:�:�ە:�`�:�:�Vn:`YR:_�5:j?:�V:x   x   ��9?�9g9��H9B~89WV39�}89�H9�g9��9w��9D��9:� :�)?:��]: �z:�:)��::ę:k�:@ę:���:��:��z:��]:�)?:�� ::��9x   x   m�w9�q;9.�9��8�S�8GU�8���8"�9wp;9Ԍw9ꤣ9���9�	:R&:�F:�&f:QT�:�:5l�:bę:ř:�k�:��:zT�:)%f:��F:S&:�	:[��9-��9x   x   �9�_�8�|8p9/8�81@/8�{8^�8ږ9tY_9D��9�!�9w�	:/}*:�wK:��j:���:=�:d��:�ݕ:���:��:a��:�j:IyK:|*:��	:!"�9� �9&[_9x   x   �[f8�R7>c�4طLط�c�"�R7jTf8���8�uM9�8�9[��9 I:2�,:['M:��j:�U�:e�:ec�:[c�:��:�U�:�j:3&M:v�,:�J:���9�7�9gtM9C��8x   x   d�׷Q�z�����;!��������z�`�׷���7R�8/�A9��9��9��:V�,:zK:Y'f:'�z:�:!�:�:�z:�'f:�zK:�,:��:k�9n �9��A9��8���7x   x   �ȸ՝�����4��@�����ȸ5�a��f�62��8��;9�e�9U�9K:F}*:˦F:��]:�[n:*�v:K�v:�\n:��]:v�F:X}*:�J:~�9�f�9��;9k��8JK�6гa�x   x   4� �4���:�o�4�Ұ �Y���'ؔ�e�����8E�;9E�9���9Z�	:T&:-?:�_R:��^:Яb:E�^:^R:F-?:U&:��	:߰�9��9��;9���8gV���ٔ� ���x   x   !UO��1\��0\��TO�c�4���
��֠�	s�����8��A9B9�9)!�9�
:z� :��5:;�D:�L:��L:��D:j�5:� :�
:8"�9T6�9C�A9;��8�����Ӡ�,�
�`�4�x   x   �Np�q�v��Np�	�\�<�;�C�
��┸=��6���8�jM96��9K��9G :dA:�S+:n6:��9:�6:<S+:B:$ :#��9���9OnM9��8A}�6r㔸��
��;��\�x   x   ����v���\�H�4�������a�i��7���8jQ_9��9��9X:p�:�� :�':S�':� :{�:�W:N��9J��9rR_9���8g��7��a�������4���\���v�x   x   �h��������ʸ�"p��I�zna8)� 9f�O9Nސ9�[�9���9�#�9��:v�:�|:h�:v�:�#�9���9�Z�9Lܐ9��O9�� 9&da8��䶢p�T�ʸ:����x   x   _��/�����<=�����qc�7�8I 9��k9��9�c�9X��9�,�9L�:��:��:��:�*�9���9Qd�9�9�k9	L 9g��8�7c��_G��-�⸟��~��x   x   ���2��𽩸��4����6��{8z_ 9�PF9F�9|��9ť�9���9���9(p:æ:p:K��9��9h��99��9�9UNF95^ 9B�{8���6Ѥ4�ѱ����⸱��[��x   x   T�ʸ%G���4�~�ٵ��J8�`�8�.9�q9��9J�9s��9GA�9�9׌:>�:x�9�?�9���9eL�9a�9G�q9�.9�_�8q�J8�H׵]�4�ZU����ʸ��Ḧ��x   x   �Jp�����%�6�J8��8�q#9	�a9�x�9�Ů9R�9W��9f�9�9n(:Ň�9�f�9��9�P�9Ʈ9�w�9��a9�s#9Z��8*|J8S��6���:p��V���[��sQ��x   x   ���/�7"�{8wW�8�o#9r�\9��9� �9�%�9���9i�9#��9�:��:��9��9���9�$�9��9s�9��\9q#9�Y�8��{8 $�7*z�R{�=.��7�Gc�x   x   �.a87�8�U 9"�.9�a9���9��9�N�9,
�9&�9A]�9G�:~�:r�:c^�9�#�9��9M�9��9P�9��a9��.9sS 9>�8Y'a8<�8ӓ7�Y[7�ʓ7��8x   x   �� 9l9 9�DF9G�q9�u�9`��9�M�9_%�9�W�9H��9:�:Z:�:%��9GW�9�%�9�O�9.��9�v�9�q9�DF9�: 9.� 9�8��8�+�8,/�8r��8��8x   x   $�O9��k9m�9�
�9�®9)$�9z	�9�W�9r��9�:y�:�
::�:y�:���9]V�9O�9C%�9®9�	�9��9��k9�O9c99�p)9!�9��9��9)q)9d99x   x   �ѐ9��9��9�D�9�N�9q��9�%�9t��9�:[	:�:۷:�Z	:��:%��9�'�9��9�O�9gE�9)��9��96ѐ9�	�9;��9�{9�%w9�,w9� {9���9V	�9x   x   iN�9Y�9��9G��9r��9k�9y]�9q:��:X�:��:g�:	�:�:�Y�9� �9��90��9��9�W�9�N�9�D�9��9���9M��9���9���9���9���9kB�9x   x   ��9���9%��9�<�9�c�9��9��:z	:�
:��:�:�
:,	:��:
��9kb�9�<�9���9���99��9k��9<��9���9�D�9o8�9�8�9{E�9��9���9r��9x   x   N�9�"�9��9P��9���9��:��:�:��:E\	:#�:�	:�:��:���9n��9\��9!�9��9�t:��:�Q	:9:c+:t�:�+:�9:�R	:a�:�s:x   x   ��:��:Wm:��:�(:�:T�::��:��:�::�::�:�(:9�:�l:N�:��::�:�l:�%:�\):��+:��+:�[):]%:�l:.�:�:x   x   ��:��:Ȥ:�:���9��9�c�9��9���9��9�^�9@��9���9�:C�:�:[�:9:9r':a�1:�::��A:��F:2(H:c�F:o�A:`�::��1:�p':�8:x   x   
x:��:o:��9�j�9`%�9�*�9�^�9�]�9%/�9J'�9Wh�9O�9�n:�:�x:��":�0:�u>:-MK:+V:w�]:X�a:��a:��]:sV:KMK:u>:k�0:9�":x   x   ��:T�:w��9�B�9���9+��9F�9�.�9T�9���9}��9�D�9V��93�:��:��":E�3:B)E:��U:Gqd:��o:�&w:s�y:�'w:�o:
qd:��U:�)E:A�3:G�":x   x   6�:�)�9\��9���9X�9�-�9�V�91Z�9�/�9,Z�9g��9b��9<*�9��:�<:��0:�*E:bY:�k:(E{:$�:��:}�:�#�:�D{:��k:�aY:*E:�0:;<:x   x   	"�97��9Ũ�95S�9�ή9��9�#�9�	�9�ͮ9oQ�9@��9���9} �9�#:w':�y>:��U:��k:�*:T�:�ы:^n�:ҋ:G�:n+:��k:\�U:�y>:�u':#:x   x   a��9�g�9T��9��9���9���9K��9W��9�9���9
f�9{��9�{:��:��1:�RK:�ud:MH{:$�:@Ѝ:;M�:M�:)Ѝ:3�:�G{:3ud:/RK:�1:`�:�z:x   x   k]�9I�9��9��q9&�a9�]9|�a9K�q9K�9��9�^�9���9�:u:ó::?V:��o:e&�:oӋ:N�:/�:N�:�Ӌ:G&�:��o:�V:m�::s:��:���9x   x   r��9�l9)_F9�.9$�#9Љ#9J�.9�aF9�l9��9<V�9� �9[	:(%:��A:��]::.w:��:�p�:�N�:�N�:�p�:��:=.w:��]:��A:b)%:`\	:��9$V�9x   x   �O9IZ 9�o 9ʈ�8a��8<��8�n 9�X 9��O9[�9��9ּ�9�C:Qg):�F:��a:�y:+�: Ջ:Eҍ:�ԋ:y�:Q�y:��a:V�F:hf):BB:���9��9?�9x   x   S� 9��8)|8��J8��J8a|8��8�� 9 �99���9+
�9�Z�9�6:	�+:Q3H:��a:b1w:�'�:��:��:(�:E0w:��a:E2H:5�+:48:�[�9�9ս�9�99x   x   ��a8G�7}�6n�͵m?�6l�7�a8�P�8`�)93F{9g�9 O�96�:��+:��F:��]:�o:VM{:s2:M{:��o::�]:��F:��+:<�:wM�9?�9�F{95�)9�S�8x   x   �}�?���f4�Of4�·�����U8���8�
 9�Lw9�ȭ9�O�9�7:ug):�A:SV:�zd:r�k:��k:�zd:�V:=�A:�g):�8:�M�9ͭ9�Mw9< 9N��8�T8x   x   ��o��0��Z����4����o���߷Ǟ�7\f�8r�9�Rw9v�9�[�9#E:�)%:��::�WK:E�U:�iY:��U:WK:ȷ::l+%:BC:7\�9��9Mw9��9�h�8!��7��߷x   x   ��ʸ��⸬��6�ʸ�4����^�\7�f�8� 9E{9y�9��9j]	:Uw:D�1:�~>:2E:1E:/>:ݗ1:�u:�]	:k��9p�9)D{9� 9�e�8��\7���T1��x   x   y�����N����>������v�7M��8��)9'��9��9�9"�:��:�y':��0:>�3:��0:�y':�:c�:6�9��9���9��)9n��8L��7����@�����x   x   ���Ć�B��Y�Ḇ8����߷�8�@�8~99��9YR�9��9;|:�&:p@:� #:�#:;@:�%:|:���9aT�9�9-x99cC�8�58��3:��<�����x   x   o�k��V�('��A���7΋8���8V�99%&|9�D�9߸�9��9�5�9>�:"/:�_:S.:A�:�6�9���9~��9�B�9�$|9��99!��8�ċ8�@�7��@��'�6�V�x   x   ��V���-������6�;8���8�%9��R9a�9�ب9'��9*��9`\�9�U:WI:"K:RT:�W�9��9~��9[ڨ9�9ϷR99!9S��8p;8�\�6��q�-��V�x   x   �8�q��̃�5<Q8\8�8EH�8Q@69��p9@S�9�:�9���9k&�9�R�9� :��:� :�U�9�*�9��9�8�9�S�9W�p9�A69xI�8�1�8,S8�m�5=���F��,�x   x   ��A�N}�6=H8Ɵ�8%��8'�%99�[9;��9�=�9�&�9���9�^�9�O�9��9�	�9VP�9�Z�9���99*�9W=�9o��9��[9Ф%9��8-��8�@8��6�VA�K����x   x   ���76�:8^/�8���8�9 9�)Q9�l�9�d�9�k�9�"�9�Q�9q��99 �9�9��9���9kT�9�"�9�j�9rc�9�m�9*Q9{7 9`��8�)�8��:8L��7�%7�}�6�W%7x   x   ζ�8$��8�:�8Ğ%9�'Q9U�9�$�9��9g�9��9=B�9n8�9)��9���9K6�9�D�9��9��9�9�#�9��9�(Q9۞%9l;�8��8���8�S8��08ߴ08V�S8x   x   g�8@9`769��[9�j�9$$�9,�9�<�9TY�9/��9b��9 ��9�C�9��9���9ϖ�9U^�9d;�9�*�9%�9�i�9�[9�56909�f�8��8��8���8m��8���8x   x   s�99%�R9!�p9V��9=b�9��93<�9Sg�9x�9bq�90��9�& :o& :��9�s�95x�94d�9�<�9��9)c�9���9��p9�R9�991�&9؜9.9�9��9��&9x   x   �|9s�9M�9q9�9�h�9��9�X�9�w�92_�9[=�9�<:RK::=:<�9�^�9�v�9�\�9��9�f�9�9�9�M�9��9w|9ͼj9T@^9��V9|RT9.�V9B^9l�j9x   x   G:�9Ш9�3�9"�9��9a��9z��9Vq�9�=�9�:�v:2v:��:,=�9s�9}��9��9�"�9�"�9�3�9�Ϩ9l9�9+��9쫔9+��9���9���9[��9ê�90��9x   x   ���9!��9.��9���9O�9�@�9$��9���9�<:8w:IB:>w:=:���93��9�C�9*R�9���9��9D��9s��9��9�ƻ9+�9-ٹ9F��9�չ9_��91ɻ9u�9x   x   t��9��9��9QZ�9+��9�7�9���9c' :	L:�v:�w:PK:�' :ՠ�9�6�9��9�W�9""�9���98��9�9.��9�_�9���9]��9���9]��9�[�9T��9n �9x   x   �*�9�S�9�L�95L�9���9q��9EE�9�' :n>:��:�=:\( :B�9���9i��9�N�9�N�9�O�9�)�9�A :5U:�\:��:��
:�5:��
:��:^:�S:�@ :x   x   ��:�Q:� :~	�9��97��9���9G��9�?�9�@�9���9���9���9��9=�9� :�Q:�:�:��:�:Un:T	!:��":F�":~	!:�m:6�:��:�:x   x   ^*:F:��:��9��99�9���9*x�9�c�9�w�9Y��9>:�9��9�	�97�:
G:i):g1:W�:�m':#'/:�N5:�>9:��::�>9:�N5:�&/:Vo':y�:.2:x   x   �[:�H:� :�P�9f��9�H�9��9~�9�|�9^��9]I�9���9�R�9N :�G:�[:Y�:"j&:�2:��<:��E:r�L:� P:��O:@�L:��E:��<:*2:�j&:�:x   x   R+:�R:�U�9�\�9�X�9���9�d�9Nk�9�c�9-��9Y�9�]�9�T�9*T:,+:N�:):�7:�E: �Q:�|[:�a:Z�c:��a:T{[:��Q:��E:!�7:�):�:x   x   O�:uV�9,�9F��9=(�9��9&C�9E�9#�94+�9���9;*�9�W�9��:?4:8l&:�7:$}H:h�W:L�d:>%n:��r:W�r:.%n:�d:��W:f{H:u�7:Cn&:4:x   x   55�9���9@��9n/�9mq�9 �9�3�9G�9lp�9�,�9#��9��9B3�9:U�:�2:i�E:��W:�"h:?�t:L�|:�]:Ɯ|:��t:�!h:[ X:,�E:82:��:h:x   x   թ�9��9B=�9�C�9Rk�9�,�9�.�9�m�9�D�9?�9���9���9�G :|�:>s':T�<:��Q:��d:��t:�:5�:~�:��:�t:o�d:m�Q:u�<:t':Z�:MF :x   x   T��9Jި9�Y�9ؾ�9�v�9��9t�9���9�Y�9�ܨ9���9�*�9\:��:�-/:w�E:��[:%)n:��|:��:�s�:��:��|:�(n:��[:]�E:�./:ي:1[:D-�9x   x   F�9#�9��p9ǜ[9�<Q94=Q9j�[9��p9�#�93G�9R(�9���9�d:,v:�V5:w�L:N�a:��r:�a:��:��:�a:��r:o�a:��L:�T5:�w:�f:���9])�9x   x   �,|9 �R9�O69��%9zJ 9�%9�L697�R9�,|9���9�ֻ9�p�9L�:!:G9:�P:��c:u�r:��|:|�:ء|:��r:��c:�P:XH9:�!:��:�n�9�ӻ9��9x   x   ��99-9[f�8���8W��8�e�8�19��993�j9���9��9���9D�
:�#:բ::�P:q�a:�+n: �t:N�t:�+n:�a:vP:��::�#:�
:���98��9U��9	�j9x   x   G��8}½8N�8�ď8�N�8ѽ�8���8p�&9p]^96��9��9��9k?:#:RH9:\�L:��[:/�d:x'h: �d:�[:L:qI9:V#:�>:C��9_�9�9�b^9��&9x   x   ֋8�7;8ȇ8�~8eC;8�Ջ8���8ж9�V9��9꺹9���9��
:^!:oX5:�F:��Q:X:5X:��Q:�F:�V5:!:p�
:q��9��9N�9��V9��9���8x   x   �|�7��6�W�5�r�6�n�7\�S8#��8]-9�nT9�	�9A�9���9`�:�w:'0/:��<:]�E:�H:��E:��<:x1/:Dy:��:f��9-�9��9�nT9�.9|»8��S8x   x   ~�@�gܸ��ĸ��@��&7�18
˳8�+90�V9v��9Ӑ�9im�9{g:#�:�w':
2:�7:I�7:�2:]w':�:�g:|o�9Δ�9���9��V9`-9���8�18�&7x   x   ��8�-��%�p����!�6%�08��8u�9[^9���9Nػ9F��9\:��:�:�q&:�
):�r&:,�:��:l\:1��9ӻ9���9o^^9��9 ��8h�08�e�6໭�x   x   ?�V�тV�S�+��ϭ��&7��S8���8��&9��j9���9�$�9Z.�9�G :o:e8:��:��:h7:�:uG :�-�9(�9���9��j9�&96��8g�S8��%7e˭�+�+�x   x   �P�7���7C@!8�}{8��8iE9Z�39%dg9�z�9c�9׏�9o��9���94�: �:o�
:+�:�:1��9���9���9K�9�y�9�bg9�39�@9��8m�{8�>!8���7x   x   ]��7�8�9T8��8a��8��9�{H9�i{9'4�9���9ob�9	T�9��9���9�:�:c��9K�9kS�9c�9���9N5�9�k{9wwH9��9���8��8{5T8>�8���7x   x   �0!8�1T8`�8Co�8�}
9K49�ob9d��9���9�|�9�O�9=��9z��9���9&��9���9���9z��9/O�9�{�9��9i��9�sb9�49E
9�s�8N�8�5T8R(!8z8x   x   !f{8��8]k�8y9K%*9�S9�P�9�h�90E�9}��9�j�9���9R0�9-��9i��9M1�9E��9�h�9ɠ�9�E�9k�9cN�9��S9#*9�w9-i�8�۝86p{8s�Z8��Z8x   x   ��8z�8�y
9G#*9�N9�Zw9x��9g�9g��9���9aH�9�A�9/��9II�9���9S@�9�K�9`��93�9�e�9���9Yw9��N9�&*9\x
9���8���8C�82_�8; �8x   x   ";9Y�9Y49?�S9 Yw9�Ǝ9ۋ�9%�9���9���9��9���9 $�9�"�9��9ǖ�9a��9p��9�9���9Ȏ9�Xw9V�S9�49V�9r69���8t��82��8�~�8x   x   ��39�qH9�gb9�M�9���9��9sC�9d@�9���9���9���9���9��9���9���9���9A��9N?�9�D�9ۊ�9A��9�O�9hb9rsH9��39�%$9k�97�9q�9�$$9x   x   �Ug9�]{9���9ye�9�d�9��9�?�9���9���9n��9�$�9I��9s��9[#�9���9ȉ�9���9?�96�9me�9Ce�9��9]{9�Qg9�X9��M9�wH9DvH9W�M9�X9x   x   �r�9Y-�9@|�9?A�9��9O��9��9n��94��9�`�92�9+��9�2�9�_�9���9}��90��9<��9��9B�9�{�9�-�98t�90��9q��9d��9˃9J��9c��9_��9x   x   nޫ9,��9�v�9M��9ҍ�9���9���9@��9�`�9���9�g�9Wf�9���9ia�9\��9��9���9���9X��9�v�9큲9xܫ9��9��9'z�9�B�9�E�9Yz�9&�9���9x   x   g��9�Z�9�I�9�f�9�E�9���9H��9�$�9n2�9Kh�9~��9Ph�91�9�#�9���9���9�H�9yd�9�J�9�Y�9;��9���9S%�9�+�9#��9���9���9�+�9�'�9^��9x   x   ���9`L�9���9ؔ�9�?�9�9��9 ��9)��9?g�9�h�9���9I��9$��9ɏ�9�=�9y��9���9�K�9���9}��97��9�D�9̈́�9�@�9�B�9��9<B�9
��9���9x   x   ��9M�9G��9-�9���9$�9��9���9w4�9���9q2�9��9�9m$�9Q��90�9���9��9��9I"�9F	 :Ss:�:��:�O:{�:�~:�t:�	 :�!�9x   x   ɐ:'��9L��9ְ�9�H�9�#�9���9�%�9�b�9d�9<&�9���9_%�9vH�9=��9���9o��9�:��:ћ:�:�:��:�^:�`:6�:;�:H:e�:�:x   x   �:&:���9D��9���9ؑ�9���9���9@��9���9���9���9c��9g��9���9>:3�:�V:VE:
:�3#:�(:t/+:�F,:.+:�(:�3#::�C:W:x   x   8�
:�:���9]1�9B�9Й�9���9Y��9?��9���9q��9�A�9P3�9I��9�:L�
:#:EV:�%:�(.:H]5:,�::�T=:sT=:2�::�^5:'.:�%::V:�":x   x   ��:ì�9W��9���9�N�9���9_��9���9��9���9�N�9���9���9V��9��:�#:�i:}�):�5:j�>:PxF:IVK:\M:}WK:6vF:��>:�5:��):=i:~#:x   x   y�:=�9t��9�k�9���9���9xE�9�E�96��9���9vk�9���9-�9͔:Y:�W:b�):�v7:��C:,�M:�UU:3+Y:�)Y:�UU:1�M:L�C:u7:��):>Y: Y:x   x   ���9�S�9~Q�9ɤ�9y��9p�9�K�9��9���9���9;S�9�S�9ԙ�9J�:�H:��%:�5:��C:��P:�Z:��`:�c:`�`:݈Z:x�P:9�C:+5:֔%:�G:w�:x   x   ���9�d�9N�9�J�95l�9���9ݒ�9n�9K�9��9�c�93��9�+�9b�:<:1,.:^�>:@�M:�Z:{yc:%h:�%h:xwc:�Z:��M: �>:v+.:Y:P�: *�9x   x   ��9���9'��9q�9� �9rЎ9��9�n�9���9`��9��9���9� :�:�8#:�a5:N|F:YU:��`:&h:��j:9&h:6�`:rXU:n{F:c5:�9#:0:� :��9x   x   ��999�9���9�T�9&hw9�iw9�X�9��9�8�9��9���9���9�y:_: (:ŕ::<[K:H/Y:�	c:�'h:/'h:�	c:�-Y:�[K:Ԗ::8(:�:�{:���9���9x   x   �|�9�t{9pb9p�S9��N9�S9~{b9#r{9��9T��9L2�93R�9��:��:B6+:/[=:M:�.Y:C�`:Jzc:��`:�.Y:�M:�Y=:Y6+:�:�:�P�9�2�9鼦9x   x   -jg9�H9�$491*9�6*9�&499�H9hgg9��9��9z9�9X��9<�:�f:N,:h[=:�]K:Y[U:J�Z:ڌZ:�ZU:�\K:�Z=:�N,:#g:��:��9�<�9y�9���9x   x   w�39��9�
9w�9�
9�9N�39�"X9���9i��9k��9�O�9�W:�h:�5+:p�::�|F:��M:,�P:z N:~F:x�::57+:qg:RV:*Q�9���9���9��9h"X9x   x   �G9���8��8��8��8�G9U9$9u�M9�̀92P�9��9�Q�9^�:"�:�(:�e5:$�>:��C:��C:��>:�e5:�(:��:��:GQ�9ћ�9�R�9:̀99�M9�7$9x   x   �8��8T/�8��8�8ȥ�80�9&�H9��9�R�9���9���9��:�:<;#:�-.: 5:bz7:m5:�..:�;#:,:��:\��9f��9kR�9��9
�H9��9���8x   x   �{8�PT8 YT8\�{8*.�8��8��9��H9�ʀ9���959�9gP�9�{:n:�:7�%:*:�*:~�%:�:�:�|:)Q�9A<�98��9k̀9�H9��9���8�(�8x   x   �L!8��8�E!8��Z8xv�8���8��9 �M9���9��94�9��9 :Ρ:�I:�[:�m:]:MJ:+�:� :0��9B2�92�9鷃9�M96�9���82��89�Z8x   x   p��7��708@�Z8�3�8[��8(3$9|X9䝈9���9k��9%��9+-�9��:�\:T':':�[:I�:,�9Y��9��9��9X��91X9�2$9`��8�"�8��Z8�58x   x   ���8�S�8���8���8�'9�x99*~`9��9�-�9�9 ��9�R�9��9���9��:ht:��:q��9`�9(S�9L��9 ��9�,�94�9�`9�s99�/9��8���8�R�8x   x   iP�8Մ�8^m�8-�
9�'9�7J9�tq9H�9��9ֹ9�Q�9�`�9N��9'2�9���9j��9�0�9��9|_�9YP�93׹9��9��90tq9�:J9��'9��
9�k�8��8�S�8x   x   I��8�i�8�u9�9A�<9��_9�C�9��9lH�9K�9k�9r;�9���9e	�9�t�9	�9���9<�9��9#�9F�9���9oD�9��_90�<9��97x9�k�88��87[�8x   x   ���8��
9Z�9Ca89W9L�y9�{�9H��9҉�9��9��9���9��9�(�9�&�9;��9{��9��9{�9;��9n��9�z�9#�y9�W9�]89M�9��
9v��8���8���8x   x   � 9Į'9��<9LW9I}u9 q�9^��9���9;s�9��9���9�_�93��9���9���9/^�9��9��9�s�9֖�9��9ho�9>u9�W9��<9��'9&"9H9�L9Ņ9x   x   �o99�0J9i�_9�y92p�9F�9%2�9� �9v��9N��9 �9N�9��9��9�L�9l �9���9&��9� �9�0�9��9�o�9�y9O�_9�-J9�l99q�-9:(9�(9��-9x   x   ds`9�kq9G@�9my�9���9~1�9 ��9�E�9H��9,N�9�S�9F�9&��9MF�9+U�9IM�9���9�D�9	��9q0�9���9�z�9�@�9�nq9�v`9��S9�nL9��I9�rL9p�S9x   x   ��9��9覗99��9���9���9SE�9���9��9h=�9]��9R��9��9��9=�9y��9��9�D�9H��9ʕ�9���9��9��9� �9��9�fw9&s9J&s9lew9ܱ9x   x   �&�9�9�C�9`��9�p�9��9���9���9���9���9���9�9g��9���98��9��9���9��9�q�9Ԇ�9�B�9�9�(�9���9@Ǔ9ct�9k��9�r�9(ȓ9���9x   x   k��9�Ϲ9`�9:�9_��9Σ�9cM�9=�9���9��9�)�9i(�9��9���9�=�9KL�9���9ʺ�9M�9��9`й9|��9��9���9��99̪9�Ϊ94��9���9��9x   x   z�9sK�9c �9A��9��9���9S�9Y��95��9*�9��9%*�9|��9���9�S�9���9���9>��9:�9K�9�z�9rz�9�1�9�p�9��9l��9s�9\p�9>3�9�y�9x   x   �J�9@Z�9�6�9H��9t]�9M�9�E�9���9��9)�9�*�9:�9���9�E�9,L�9-\�9���9�7�9 X�9AJ�9-��9_�98B�9�B�9���9���9TF�9wA�9g�9���9x   x   >�9F��9q��9%��9���9q�9���9��9���9@�9���9���9\��9��9���9ʭ�9:��9L��9��9��9���9���9�n :B:'�:�}:�m :Ĵ�9|��97��9x   x   x��9�,�9��9�&�9��9�9�G�9���9���9���9���9=G�9n�9���9`%�9$�9j,�9��9pU:�:�
:��:E�:u:x:��:_�:�
:Z:�V:x   x   ��:}�9+r�9�%�9ф�9<N�9PW�9�?�9��9e@�9bV�9uN�9S��9H&�9�s�9_~�9�:�J	:�:w3:��:S�:v2:^ :{1:!�:��:}5:��:�J	:x   x   �q:��9J�9��9[_�9��9_P�9��9���9!P�9��9q_�9���9 �9x�9�p:Q_:�:��:X�!:BM':AV+:Uo-:9o-:@W+:MN':��!:��:@�:_:x   x   ��:V.�9-��9o��9B��9>��9���9x��9���9U��9W��9��9��9�/�9?�:�_:c:Ձ:�*':R�.:��4:�o8:�9:Bp8:�4: �.:�*':�:c:�_:x   x   ���9��9=�9��9S��9i��9�I�9+J�9���9���9���9N=�9^��9z��9jL	:K�:��:W):s�2:��::C@:s;C:�:C:�C@:��::��2:�):N�:˶:�L	:x   x   �9�_�9@	�9��9�w�9��9ч�9��9Ox�9�9 	�9�^�9!�9aX:��:��:0,':?�2:8�<:�PD:x5I:L�J:\5I:�QD:?�<:*�2:-':O�:��:�W:x   x   S�9�Q�9��9:��9ߛ�9�6�9�6�9ۜ�9G��9c�9�R�9R�9���9+:�6:D�!:��.:2�::�QD:�HK:��N:'�N:GK:�QD:��::��.:ε!:�7::���9x   x   I��9�ٹ9�I�9��9���9$�9���9G��9�J�9�ع9���9,��9���9c�
::�P':��4:�E@: 7I:��N:��P:��N:�8I:�D@:��4:�Q'::��
:8��9���9x   x    ��9�9̮�9��9�u�9�v�9w��9⮗9��9௴9R��9��9ͽ�9ª:�:�Z+:�s8:�>C:��J:��N:��N:@�J:�=C:Qt8:4[+:�:Ы:V��9V�9F��9x   x   /�9F�9I�9Q�y9=�u9��y9�H�9��9 2�99��9�<�9GM�9pt :��:�7:St-:��9:�>C:Y8I:9IK:�9I:d>C:w�9:�s-:�7:A�:�r :�L�9;?�9í�9x   x   �9�{q9t�_9."W9	)W9@�_9rq9�	�9�ė97��9P|�9�N�9D�:u:+
 :�t-:)u8:�G@:iUD:TD:�F@:]u8:�s-:�
 :�:˅:�O�9�{�9i��9�Ɨ9x   x   ��`9wBJ9��<9^i89��<9�<J9a�`9&�9aѓ9�ū9|%�9���9c�:�:�7:�\+:0�4:�::ۙ<:T�::�4:v\+:w8:�:Q�:$��9q$�9�ū9ғ9��9x   x   �y99�'9��9T�9N�'96{99>T9yw9�~�9>ת99
�9���9�:��:5�:�S':7�.:�2:Ƨ2:��.:�S':V�:��:�:>��9��9�٪9&�9�uw9AT9x   x   59��
9��9��
9>.9t�-9�~L9u8s9_��9y٪9"�9lR�9�s :x�:�:"�!:�/':):d0':R�!:�:�:'s :UP�9X$�9R٪9!��9;s9�L9��-9x   x   _��8	w�8�z�8%��8j�9Z%(9��I9d7s9w|�9�ƫ9j{�9�L�9c��9��
:�::�:E�:�:*:�9:��
:���9M�9�{�99ū9�~�95:s9��I9�#(9]�9x   x   [��8��8���8��8�V9�(9��L9Juw9�Г92��9�=�9��9��9:��:��:�f:ǹ:0�:�:���9��9�>�9a��9�Г9	sw9�~L9�"(9�]9�8x   x   V�8�Y�8e�8Q �8D�9T�-9�T9%�9�9¬�9*��9���9z��9[:�N	:�b:�b:�N	:>Y:���9���9���9O��9�ė9��9(T9�-9��9Z�8�h�8x   x   Y49��9�� 9B19��G9wd9b~�9���9��9Or�9}4�9=�9���9ƴ�9'��9@� :D��9���9���9r=�9�4�9�s�9��9J��9�}�9�d9G�G9�D19&� 9_�9x   x   "�9� 9��)9d�<9��T9��q9qo�9�#�9�q�9nr�9�H�9��9��9H^�9���9��9_�9��9��9H�9�q�9�p�9b$�9�p�9��q9��T9��<9,�)9�$9�9x   x   �� 9t�)9��89 UM9)�f9�9t��9��9��9N>�9��9�~�9u��9��9��9���9r��9~�9��9|?�9j�9�9���9��9�f9yVM9��89��)9+� 9�9x   x   �=19d�<9�SM9�b9�C|9�~�9o�9�ë9)<�9G��9�]�9
��9N��9�c�9�c�9ǳ�9���9�]�9��9n;�9�ë9��9��9dB|9v�b9�QM9�<9�@19��+9n�+9x   x   ��G9�T9!�f9B|9���9�h�9�ݦ9WM�9�"�9.��92�9+�9)�9���9��9+�9�1�9��9�$�9�L�9Qݦ9kg�9���9�C|9ɉf9`�T9'�G9 @9�w=9N@9x   x   �d9��q9��9U}�9�g�9�B�9�Z�9wA�9;�9���9T-�9�9��9J�9��9J-�9��9�9�9�@�9�Z�9�C�9)h�9�}�9��9/�q9d9E�Z9n�U9�U9
�Z9x   x   �y�9�k�9���9X�9:ܦ9Z�9q�9j�9��9��9~�9��9
v�9��9��9ŕ�9��9�9�9:Y�9)ܦ9D�9���9�l�99z�96�z9y�t9x�r9�t9d�z9x   x   Q��9�9B�9���9�K�9i@�9��9C�9�f�9���9��92��9[��9���9���9ye�9�C�9E�9@�9�K�9���9��9��9��9��9V�9ܣ�9(��9{W�9J��9x   x   ��9�l�9�9'9�9� �9�9�9G�9�f�9���9GR�9�M�9�D�9�N�9�R�9���9ef�9��9l9�9<!�9�8�9��9<m�9��9���9�u�9N��9��9q��9�t�9��9x   x   l�9$m�9:�9��9���9#��9Y��9L��9AR�9Im�9��9��9<l�9�P�9U��9ǔ�9���9"��9X��9�9�9ll�9�k�9�1�9F�9�Y�9Δ�9#��9[�9~�91�9x   x   �-�9�C�9��9�Z�9�/�9,�9� �9���9N�9��96��9��9�P�9���9� �9	,�9[/�9~Z�9�99D�9�-�9ӡ�9m��9��9���9���9 ��9~�94��9B��9x   x   z6�9I�9`z�9!��9:)�9�9f�9h��9ME�9'	�9@	�9{C�9���9#�9�
�9*)�9��97z�9��9y6�9o��9:��9���9���9���9���9ˌ�9���9���9���9x   x   U��9h �9���9ɰ�9��9d�9Dv�9��9�O�95m�9zQ�9.��9bv�90�9K�9j��9���9��9n��9��9��9f+�9��9�U�9���9�U�96��9b+�9��9(��9x   x   ��9�Y�9���9�a�9���9y�9��9U��9AT�9,R�9&��9=�9��9���9�a�9���9�Y�93��9���9�B:�:�x:�5	:$
:�#
:"6	:iy:@:AB:��9x   x   ��9ܧ�9���9_b�9��9��9Z�9���9Ǟ�9���9��9��9��9=b�9g��9ק�9V��9:8�:��:�:�{:\[::�[:"{:�:5�:Q�:{:x   x   � :���9T��9{��9�+�9�.�9��9Ph�9oi�9ӗ�9�.�9�+�9���96��9���9�� :ؕ:�r:�9:v:��:!�:D� :4� :N�:�:�t:�9:�s:��:x   x   ��9]�9���9C��9\3�9���9	�9|G�9W�9���9&3�9���9���9k\�99��9Z�:��:|:[�:��!:�W&:xD):	G*:�C):�W&:��!:��:�:m�:��:x   x   p��9��9R~�9k_�9���9'=�9��9��9�=�9ݦ�9 _�9�~�9��9ٰ�9�:�s::�Q:L�$:�*:�_/:�1:ګ1:w`/:��*:��$:SR:1:�s:�:x   x   w��9��9��9e��9�'�9�D�9��9E�9�&�9��9��9s�9���9���9L�:�;:��:��$:a�,:f�2:�U6:�7:%T6:.�2:P�,:M�$:��:�;:��:Ҍ�9x   x   S=�9I�9�A�9�>�9�P�9�_�9�^�9�Q�9?�9#@�9�J�9�<�9a��9�E:��:Ux:��!:Y�*:�2:��7:n�::��::��7:2�2:��*:��!:	x:-�:�E:���9x   x   j5�9�s�9A�9uǫ9��9�H�9�9=ǫ9R�9�s�9F5�9���9!�9@:1�:��:(Z&:�a/:�V6:�::�7<:$�::wW6:2a/:Z&:��:��::< �9��9x   x   ?u�90s�9t�9�9}l�9�m�9��9��9�t�9�s�9��9v��9�3�9�|:�:��:|G):��1:ȥ7:��::��::�7:��1:�G):�:�:�|:�4�9e��9E��9x   x   ���9J'�9� �9���9Z��9���9��9"&�9���9�9�9$��9���9��9_:	:�_:;� :�J*:ˮ1:xV6:B�7:�X6:r�1:�I*:H� :�_:�:	:��9���92��9�8�9x   x   ���9�s�9��9�K|9�N|9�9�s�9���90��9�9!�9���9S_�9�(
:�:}� :�G):�c/:ڎ2:7�2:�b/:�H):�� :�:^(
:�_�9��9��9��9⚣9x   x   ��9�q9�f9��b9ٔf9��q9?��9?��9	~�9�b�9{��9��9���9�(
:�`:��:[&:5 +:#�,:�+:�[&:�:h`:�(
:\��9^�9��9�b�9�}�9Q��9x   x   `d9��T91^M9�ZM94�T9j"d9�z9�]�9Ř�9睳9*��9��9�_�9!;	:�:��:��!:l�$:�$:��!:d�:��:;	:+`�9y�9D��9���9���9'^�9F�z9x   x   ��G9H�<9��89��<9w�G92�Z9��t9j��9���9��9���9���9"��9E~:��:y:r�:�U:0�:�y:\�:�}:���9W��9���9���9s��9���9�t9\�Z9x   x   H19�)9��)9�H19�@9u�U9B�r9Y��9d��9�c�9� �9&��9�4�9�:��:�=:C
::�=:��::�5�9��9x�9Kb�9u��9E��9��r9Q�U9m@9x   x   �� 9�(9�� 9�+9p�=9<�U9��t9"^�9|�9��9���9)��9�"�9cF:+�:4w:^�:Yv:`�:G:�!�9���9��9��9�|�9]�9n�t9i�U9��=9��+9x   x   ��9ѯ9A�9.�+9�@9�Z9��z9U��94��9J8�9ȩ�9_��9���93��9�:��:ژ:�:8��9���9O��9���9j7�9]��9���9�z9u�Z9R@9��+9i�9x   x   !�B9��E9�SN9oi\9��o9o��9k^�9~�9:q�9
|�9)��9{��9D��9��9E�9#�9
F�9x��9֫�9���9?��9\~�9r�9,~�9]�9ǜ�9�o9�i\9gRN9��E9x   x   ��E9�%K9�
V9:�e98?z9�L�9���9���9�մ9ح�9 ��9p��9`�9�>�9���9t��9�@�9a�9ܣ�9���9۫�9�Ӵ9���9���99M�9�Az9��e9�	V9\(K9q�E9x   x   .QN9�	V9�b9C�s9�e�9Ȍ�9���9���9N�9�v�9���9���9��9 X�99�9X�9���9���97��9�v�9��9��9x�92��9|d�97�s9��b9�V9�ON9�K9x   x   �e\9��e9�s9�Ȃ9�\�9pG�9�
�9Q�9�ٿ9���9��9�p�9�9�98�9:�9&9�9�q�9��9���9�ٿ9�9�
�9�H�9[^�9�Ȃ9)�s9<�e9f\9GxW9�vW9x   x   q|o9V;z9�d�9S\�9���9��9��9=к9 $�9�V�9���9g�9&y�9g��9�w�9�h�9��9�V�9-%�9�Ϻ9}�9��9���9�[�9he�9�:z9@~o96�h9
�f9��h9x   x   1��9�I�9ڊ�96F�97�9(��9�A�9���9�{�9��9I��9���9,$�9z$�9 ��9>��9��9�z�9y��9aB�9��9��9�G�9���9sJ�9n��9&c9�w{9 y{9-f9x   x   �Z�9���93�9��9��9VA�9С�9C��9H��9y��9=��9��9��99�9���9��9`��9���9E��9�A�9��9)�9��9���9�Y�9.�9���9�Ӊ9�9Y-�9x   x   �y�9൥9��9�9�κ9���9��9���9�p�9��9�Z�9o=�9�<�9�[�9���9o�9���9Ȕ�9��9Ϻ9��9��9ڵ�9ez�9�u�9��9tY�9�Z�9���9�u�9x   x   Ul�9�Ѵ9��93׿9U"�9|z�9���9up�9/F�9��9b�901�9|a�97�9jG�9�p�9n��9{�9V!�9�ֿ9� �9�д9�k�9��9rk�9��9�a�9�ߨ9�j�9��9x   x   �v�9u��9Js�9��9�T�9l�9ə�9Ǥ�9��9jr�9 ��9]��9uq�9g�9���9V��9Q�9gT�9���9�q�9���9�x�9q��9-�9ݺ9ZE�9nE�92ݺ9��9���9x   x   ���9��9$��93�9���9&��9���9Z�9%b�9��98+�9.��9(d�9�Z�9���9L��9���9��9ޒ�9���9Q��9z��9e��9���9YL�9{=�9M�9��9���9x��9x   x   ��9��9��9!n�9qe�9���9��9�=�9�1�9���9q��9J0�9�<�9��9)��9�f�9�p�9���9��9t��9�u�9�:�9��9A��9��9��9���9��9E;�9�u�9x   x   ��9�[�9Ð�9�7�9�w�9�#�9��99=�9-b�9=r�9�d�9=�9��93#�9{w�9�5�9׎�9^�9ܥ�9vG�90��9�\�9�`�9���9��9l��9_`�9}\�9���9�F�9x   x   =��9�:�9lU�9b6�9���9u$�9��9�\�9m�9��9�[�9��9�#�9���9�7�9
X�9�:�9��9�e�97�9�W :�B:��:�X:�W:S�:�B:=W :o8�9�e�9x   x   �@�9���9��99�9�w�9���9���9;��95I�9z��9=��9���9�x�9?8�9���9|��9�@�9?=�9{.:�:��	:��:fN:��:"O:��:��	:��:.:�;�9x   x   ��9���9�V�9�8�9i�9���9���99q�9
s�9Ҝ�9���9�h�9s7�9aY�96��9� �9�:W:��
:�:w�:�:d8:�8:��:�:�:��
:6X:I�:x   x   QC�92?�9��9r�9=��9�
�9���9���9���9��9���9�s�9a��9�<�9DB�9~�:ul:A*:��:�1:s�:h:��:>:��:Y2:܍:):�k:̢:x   x   ���9�`�9���9��9�X�9Z}�9���9H��9�~�9BX�9��96��9qa�9��9�?�9�W:�*:��:7�:�u:��!:+�#:��#:u�!:�t:՝:<�:6+:X:?�9x   x   ۪�9��92��9n��9�'�9���9��9&��9�%�9��9n��9���9��9�i�9*0:�
:��:��:��:�e$:�V':�X(:�U':�e$:&�:�:�:1�
:�/:�k�9x   x   ���9|��9xx�9ܿ99Ӻ9=F�9�E�9�Ӻ9�ۿ9w�9���9���9�L�9�;�9�:�:p3:�v:Ef$:��(:l�*:��*:�(:�e$:Dv:I4:�:�:�:�9�K�9x   x   ���9S��9�90�99�9o��9j�9��9��9ϭ�9M��9�{�9��9UZ :2�	:ˆ:e�:~�!:�W':��*:��+:��*:kW':��!:��:m�:��	:f[ :���9@{�9x   x   ��9�մ9���9�9��9��9n�9���9	״9>�9��9�A�9Jc�9�E:��:��:�: �#:&Z(:��*:L�*:�Y(:�#:�:�:��:E:5a�9%C�9��9x   x   �s�9���9���9aL�9�9�L�9Y��9���9"r�9]��9��9	�9�g�9D�:�Q:�;:S�:ԩ#:fW':+�(:;X':t�#:��:F<:�Q:J�:^j�9	�9��9���9x   x   ��9g�9q��9Pb�9�`�9؎�9n �9���9��9o�9"��9��9Ů�9�\:'�:(<:B:�!:�g$:g$:��!:y:�<:��:/\:\��9ܫ�9���9�9��9x   x   _�9�O�9�g�9�̂9j�9�O�9s_�9@|�9mr�9��9 T�9��9�%�9�[:�R:B�:��:Pw:\�:�w:��:��:<R:Y\:�(�9�
�9�T�9p�9�q�9s|�9x   x   ���9�Fz9��s9�s9�Cz9���9�3�9���9��9�L�9WE�9�9���9R�:��:h�:}5:��:E�:�5:��:��:��:���9�
�9�E�9OL�9��9���9�4�9x   x   ��o9J�e9��b9��e9҆o9+m9���9�_�9^h�9�L�9�T�9���9\h�9�F:��	:C:ސ:��:�:S:
�	:�E:
k�9��9�T�9-L�9�i�9`�9r��9wn9x   x   �l\9V9 V9�l\9>�h96�{9Dى9�`�9�9?�9q��9Y
�9d�9�Z :6�:��
:<,:|-:��
:e�:=\ :b�9H	�9s��9	�9^�9�_�9'ډ9��{9,�h9x   x   �TN9�+K9*TN9*~W9Y�f9ȁ{9맊9-��9�p�9<�9��9IB�9���9?�9'1:�Z:n:�Y:O1:`<�9���9lC�9r�9o�9q�9���9§�9.�{9Ϭf9�~W9x   x   �E9��E9q�K9�{W9%�h9�m9�1�9�z�9u�9���9���9�{�9�L�9�k�9A�9��:��:�A�9�m�9�L�9�{�9���9���9��9{�9Q3�9l9c�h9�}W9��K9x   x   �zj95�l9�t9��9���9S�9U�9�9�$�9]�9��9i}�9�$�9xl�9L��9�{�9���9�h�9n$�9m{�9I�9�_�9M%�9�9.T�9V�9���9h�9Zt97�l9x   x   >�l9�q9�z97�9yp�91��9���9A.�9I��9���9�=�9<-�9	�9���9`��9���9���9W �9�-�9]@�9��9���94-�9���9O��9Qr�9C�9��z9�q9�l9x   x   �t9��z9���9ƭ�9"y�9���9��9k?�9�ؾ9���9���90+�9y�9]r�9%��9�r�9�w�9`*�9"��9H��9^ھ9�A�97��9?��9�v�9x��9D��9�~z9Ht9��q9x   x   h�9�97��9��9��9���9DA�9% �9{�9k.�9���9��9rC�9���9̲�9�A�9��9w��9
/�9�|�9���9G@�96��9��9��9���9�9\�9;�{9!�{9x   x   ���9�n�9x�9@�9Re�9׼�9Ps�9f/�9!m�9���9G��9��9$f�9��9 d�9��9���9���9�k�9l/�93v�9ν�9\c�9T�9�w�9�l�9	��9�E�9dW�9hC�9x   x   ��9��9a��9���9S��9�M�9��9Ԓ�9���9
r�9���9��9���9#��95��9���99t�9��9��9��9 J�9#��9��9՚�9/��9��9��9��9y�9v��9x   x   �Q�9��9���9�?�9`r�9h�9��9���9w�9��9�-�9,��9p��9���9�,�9���9�s�9���9��9j�9t�9,=�9��9��9�P�99�9R��9,+�9���9S�9x   x   X�9-+�9�<�9@��9.�9��9\��9���9k��9�,�9��9���9��9 �9�,�9���9���9k��9��9�-�9���9>�9�+�9��9n��9yt�9^N�9N�9�s�9���9x   x   z �9ܧ�9�վ9�x�9�k�9���9{v�9-��9���9���9��9�@�9��9	��9	��9��9lt�9φ�9�i�9�x�9�׾9���9f �9�U�9�G�9��9ם�9|�9aI�9�T�9x   x   �X�99��9���9#,�9R��9 q�9���9],�9���9���9���9��9?��9���9�+�9n��9Cs�97��9v/�9���9Y��9�[�9]�9���9�ݿ9�_�9�^�9ܿ9���9)_�9x   x   ��9�9�9~��9���9���9���9q-�9��9��9���9��9���9��9��9i.�9s��9-��9��9���9�<�9��9� �9��9�)�9���9��9���9�*�9R��9�!�9x   x   �x�9�)�9M(�9�}�9l�9G��9���9���9(A�9$��9ݑ�9�B�9e��9>��9���9��9f��9=(�9,*�9@w�9���9!��9�=�9���9��9��9���9@�9��9��9x   x   c �9��9^v�9�A�9e�9��9l��9<��9u��9ޚ�9q��9���9���9��9�d�9�>�9)t�9 �9��9c6�9i�9vc�9���9^��9�Q�9>��9���9�c�9�j�9�3�9x   x   �h�9e��9p�9���9;��9��95��9��9���9���9f�9���9f��9���9���9�s�9��9h�9N�9(1�9~��9h��9��9��9��9��9��9~��903�9KM�9x   x   ���9ĕ�9`��9ձ�9�c�9���9y-�9�-�9z��9�,�9�/�93��9�e�9'��9f��9A��9���96��9e]�91b:w�:L�:��:�:��:��:b�:�`:s^�9~��9x   x   �x�9���9�q�9�A�99�9���9��9_��9���9n��9d��9f�9�?�9�t�9Ԕ�9Bz�9G��9�@:��:�,:��
:9�:@�:A�:+�:�
:�-:�:�@:2��9x   x   ���9J��9Lw�96��9���9�u�9�u�9���9�v�9�u�9���9Ƃ�9Bv�9ױ�9#��9���9�":��:u�
:�:Aq:;:��:�9:�r:��:�
:P�:�":f��9x   x   *g�9��9t*�9N��9(��9���9e��9@��9މ�9X��9/��99+�9��9�j�9)��9�A:��:��:��:tX:::p:4q:�:@X:Ɛ:�:��:A:���9x   x   �#�9�-�9���9{0�9�m�9���9���9z��9ym�923�9E��9�-�9F"�90Q�9`�9��::�
:�:,V:��:�P:E:�P:$�:�V:�:X�
:��:�a�9�S�9x   x   O{�9�@�9���9�~�9�1�9�9��9�1�9�|�9��9A�9�{�9�:�95�9�c:.:5�:@Y:) :�K:��:��:�L:B :vX:�:�.:c:j1�9�9�9x   x   ��9)��9/ܾ9O��97y�9�M�9�w�9!�9,ܾ91��9}�9z��9�m�9��9��:n�
:�r:f	:rQ:M :%�:! :,P:
:�r:��
:H�:y��9p�9���9x   x   �`�96��9�C�9C�98��9«9zA�9�B�9���9�`�9
&�9���9�h�9���9��:j�:�<:�q:k:��:} ::Xr:\<:H�:ъ:$��9�e�9n��9�%�9x   x   �&�9+/�9²�9L��9g�9Cã9��9�0�9�%�9�b�9��9�C�9���9���9a�:��:��:�r:R:�M:�P:�r:"�:��:��:5��9R��9�C�9��9�b�9x   x   ��9���992�9"�9%��9���9�9C[�9���9�/�9+��9���9��9�:��:<:�	:� :|:�
:�<:��:*:��9��9���9�/�9���9�Z�9x   x   �U�9���9Sy�9�9�{�9���9~U�9˭�9�M�9��9���9A�9CX�9,�9��:��:fu:^Z:~X:�Y:�s:��:�:��9�Z�9t�9�9f�91M�9��9x   x   ��9tt�9#��9հ�9op�9P�9��9�y�9V�9�e�9{��9M�9���9x��9��:��
:�:�:��:X�:��
:n�:���9`��9��9l��9)e�9c�9�y�9^��9x   x   d��9D�9ȉ�9��9���9-��9�9�S�9���9�d�9K�9!��9N��9C��9V�:t0:u�
:�:��
:�/:!�:2��9���9��9�9e�9���9�R�9��9���9x   x   ��9_�z9�z9�9%I�9x�9�/�9S�9��9��9�0�9:F�9�i�9\��9�c:��:x�:P�:R�:�d:���9mf�9�C�9s/�9�9�9�R�9m0�9��9�I�9x   x   t9��q9t96�{9nZ�9�9��9Px�9xN�9
��9���9���99p�9�8�9nc�9�B:�$:�B:*d�9�2�9�p�9���9͋�9��9�L�9y�9�9J�9NY�9��{9x   x   ,�l9�l9��q9P�{9F�9���9��9묦91Y�9d�9�&�9*��9�8�9�Q�9å�9���9t��9��9wU�9d:�9���9?%�9�a�9�Y�9�9A��9���9-I�9�{9�q9x   x   ���9G��9l��9X��9�M�9(��9Y"�9!��9�g�9�O�9���9H�9b��9���9��9��9��9K��9���9��9��9�Q�9/h�9���9"�9���90J�9i��9��9:��9x   x   Ֆ�9��9�R�9�ޑ9!��9~n�9��9h��9�F�9K�9L��9S��9�D�9���9��9��9���9_F�9���9��9�I�9�E�9K��9��9m�9���9��9�T�9k��9���9x   x   ���9]R�9e��9���9���9c�9Ń�9��9*��9��9q��9���9���9��9��9j�9@��9���9���9h��9���9��9���9�c�9��9���9\��9�P�9t��9T��9x   x   ���9�ݑ9 ��9P˜9��9W6�9��9��9�V�9&O�9,<�9���9���9Ӧ�9���9^��9]��9�<�9iP�9�X�9��9��9:5�9��9˜9���9��9���9��9��9x   x   &L�9���9��9�9��99ɲ9lȺ9)��9iS�9��9��9�%�9���9��9���9N'�9^��9�9Q�9���9�ɺ9�ʲ9��9j�9��9J��9�J�9��9�C�9��9x   x   ���9�l�9�a�9n5�9�Ȳ9�ѹ9���9���9�^�9��9���9���9�B�9D�9��9���9���9`�9���9W��9�ι9Cɲ9�6�9�a�9�n�9[��9��9���9���9Q�9x   x   ��9[�9���9��9�Ǻ92��9��9���9D�9��9~�9k0�9���9�.�9��92��9�?�9V��9�9F��9�ɺ9x�9��9��9��91V�9���9
�9[��9pV�9x   x   ��9���9��9z��9��9��9:��9���9X��9�*�9���9���9w��9��9[*�9���91��9���94��9z��92��9�9���9q��9�ծ9o�9`�9��9��9;֮9x   x   Ld�9�C�9ڑ�9�T�9$R�9�]�9�C�9&��9��9~,�9��9��9��9$,�9���9���9"A�9�^�9cQ�9*U�9��9<A�9�c�9r�95r�9]y�9�%�9�{�9�s�9�9x   x   CL�9H�9���9@M�9R�9$��9p��9�*�9m,�9N��9�Z�9$[�9��9�.�9�(�9í�9���91�9RP�9ĥ�90H�9EO�9{��9�{�9#��9�K�9�I�98��9�{�9*��9x   x   K��95��9���9G:�9���9���9��9f��9��9�Z�9���9�Z�9Ƥ�9��9��9�9;��9:�9���9o��9���9���9�}�9;�9��9��9S�9";�9�|�91��9x   x   ��9M��9���9ӽ�9x$�9���90�9���9��9[[�9�Z�9b�9Y��9�-�98��9$%�9��9k��9���98�9�9��9���9Y��9D�9��9���9��9|��9�}�9x   x   ���9�A�9���9��9���9GB�9���9���9���9[��91��9���9`��9C�9_��9 ��9��9�B�9���9���9!d�9_��9;�9f�9 Z�9��9F:�9���9�f�9���9x   x   ���9(��9�9���9u��9�C�9/�9��9�,�9�/�9���9d.�9YC�9��9w��9��9���9��9��9D*�9��9�l�9{$�9��9j�9%�9�l�9
�9{+�9�9x   x   ��9��9l�9���9d��9"��9>�9M+�9���9�)�9��92��9#��9ާ�9��9��97��9,-�9\��9J�9���9a :HI:��:�H:%a :���9��9���9�-�9x   x   ���9��9k�9���9�'�9-��9J��9��9��9]��9R��9�&�97��9]�9f�93��9��9-��9���9g�:��:(:��:��:�(:��:݁:W��9v��9��9x   x   B��9���9���9���9��9���9*A�9	��9"C�9���9R��9���9���9,��9<��9���9H�9\Y:/�:V�:F�	:�@:��:�?:��	:��:��:�Y:gI�9���9x   x   ��9�E�9���9[=�9;�9�a�9Y��9��9a�9��9�<�9٪�9�D�9���9�.�9N��9�Y:�{:n.	:�/:I:�b:�c:zH:M0:�.	:�{:�Y:^��9\-�9x   x   ��9���98��9�Q�9�R�9���9x�9���9OT�9`S�9���9���9q��9	�9���9h��9ɽ:�.	:��:��:&�:GJ:S�:�:��:/	:(�:��9���9�
�9x   x   ��9v��9|��9xZ�9���9���9-��9���9�X�9G��9���9�	�9_��9l-�9 �9��:B�:W0:9�:�v:r�:<�:�w:��:�/:��:f�:��9
)�9��9x   x   B��9�J�9q��9"��9`̺9cѹ9ͺ9���9���9L�9���9��9h�9y�9���9w�:��	:J:Ư:��:��:��:ۭ:�J:��	:��:p��9�9�i�9��9x   x   �R�9G�9��9��9LͲ9v̲9
�9�9`E�9�S�9T��9w�9���96q�9c :�):{B:�c:-K:��:��:qL:wd:eA:[*:�c :�n�9t��9E�9Z��9x   x   8i�9���9���9�7�9��9�9�9Ⅿ9��9Gh�9��9���9|��9�?�9)�9tK:��:<�:+e:p�:�x:W�:�d:�:��:8J:*�9gB�9���9?��9ȫ�9x   x   ߍ�9g�9�e�9L�9��91e�9��9Ǝ�9$�9�9@�9w��9��9�
�9�:��:�A:J:_�:��:�K:�A:��:ƙ:��9D�9���9�>�9��9�#�9x   x   o#�9�n�9Q��9�͜9���9<r�9#�9�ٮ9�v�90��9��9�#�9I_�9�
�9K:�*:|�	:�1:��:�0:r�	:�*:vJ:��9�_�9�#�9��9���9Jv�9?ۮ9x   x   䗝9M��9ï�9D��9h��9���96Z�9��9&~�9�P�9�9"�9=�96*�9�c :ʥ:{�:�0	:u0	:��:a�:cd :�*�9|�9�#�9��9nP�9��9n�9�X�9x   x   kK�90�9q��9 �9N�9���9���9�"�9�*�9�N�9u�9���9}?�9�q�9H��9�:u�:*}:p�:[�:���9�o�9�B�9��9��9]P�9�)�9�!�9��9���9x   x   i��9UV�9�R�9搎9��9Ԡ�9��9!�9���9��9@�9���9���9��9
�9Y��9N[:t[:X��9a �9#�9��9��9n>�9Q��9��9_!�9��9���9��9x   x   Ǡ�9���9��9��9rF�9���9إ�9�	�9�w�9`��9A��9( �95k�9�/�9���9	��9jL�9���9���9@*�9�j�9|�9��9���9�u�9��9
��9j��9vF�9L�9x   x   ���9W��9���9D�9��9 ��9�Y�9�ٮ9�!�96��9_��9���9ѧ�9��91�9���9��96/�96�9���9A��9��94��9-#�9Lڮ9�W�9��9�
�9��9���9x   x   � �9��9pv�91��9g<�9e�9-��9U��9��9���9"�9q��9X�9$��9���9��9���9��9��9̱�9��9x��9Д�9(��9���9P�9�9�9���9�t�9h�9x   x   .�9���9P��9lS�9�E�9FA�9��9�d�9���9�!�9{��9�c�9���9�l�9�W�9�T�9Ol�9���9�e�9���9]!�9p��9�d�9��95>�9E�9�U�9��9S��9u�9x   x   �u�9ഘ9�R�9�K�9�]�9JL�9*ߵ9v½9���9`�9e��9�E�9�~�9��9��9:�9�}�9�C�9ڬ�9��9���94ý9Gݵ9�L�9�_�9�K�9PO�9���9}v�9���9x   x   ��9�R�9 K�9�i�9�i�9��9TE�9���9���9:�9[��9|L�9up�9��9v�9fo�9pN�9��9�9u��9���9�F�9<�9j�9�g�9aL�9�V�9Q��9�3�9n4�9x   x   �:�9�D�9�\�9�i�9�;�9a~�9w�9+��9��9K�9���9Ko�9K��9Mi�9s��9p�9N��9 J�9���9)��9-�9h�9�;�9�i�9�^�9eA�9�8�9<Z�9��9vX�9x   x   ��9�?�9%K�98�9~�9X.�9��9d��9d��9���9b4�9���9��9Y�9���9�2�9Ί�9���9k��9��9-�9j}�9��9�J�9�?�9��9��9�ˣ9]ͣ9E�9x   x   ���9��9�ݵ9BD�9��9l�9��9��9N�9a��9=f�9e�9��9��9-g�9C��9��9���9�
�9��9S�9�C�9�ݵ9��9���9m��9�F�9 Ӫ9^F�9m��9x   x   ˖�9�b�9���9���9C��9ݳ�9���9��9W��9��9�y�9�h�9�j�90{�9���9���9q��9���9���9ŉ�9���9���9Xd�9���9Zj�9�9�1�981�9��9k�9x   x   &��9!��9���94��9׽�9���9��9,��9�J�9c(�9ET�9^��9|R�9�'�9CK�9���9��9/��97��9n��9w��9���9T��9��9lg�9+��9�E�9⓼96f�9���9x   x   ̄�9l�9L�9��9�I�9ɇ�9��9ܖ�9K(�9�?�9g��9���9lA�9�)�9���9F��9��9�G�9��9� �9 �9��9;�9s@�9	��9xA�9>�9Ӕ�9B�9u:�9x   x   ��9���9J��9»�9���9�3�9�e�9�y�9<T�9k��9��9��9Q�9�{�9gg�9�1�9n��9n��9ê�9���9��9�x�95 �9���9'��9���9}��9W��9&�9�y�9x   x   s��9,a�9�C�9�J�9Dn�9��9�9�h�9v��9��99��91��9[i�9,�9���9o�9�K�9qB�9hb�9ΰ�9E�9M��9���92:�9Ge�9Ge�9�8�9���9���9@�9x   x   ��9A��9}�9'o�9n��98�9��9�j�9�R�9�A�9lQ�9�i�9J��9��9���9�l�9y}�9��9G�9��9[��9�A�9G>�9���9��9U��9!?�9M?�9���9I��9x   x   |��9�j�9R�9��9�h�9%�9��9�{�9?(�9G*�9(|�9��9��9�e�9��9��9�i�9��9��9��96]�9'J�9��9�V�9?W�9"��9bJ�9^�9��9���9x   x   ���9�U�9=�9��9;��9���9�g�9z��9"L�9w��9Oh�9|��99��9��9 �9�T�9��9O��9�u�9���9i��9c-�9��9�%�9���9,�9���9��9kx�9b��9x   x   5��9SS�9a�9o�9#p�9<3�9��9���9���9���9�2�9=p�9�m�9��9 U�9B��9x��9���9�z�9O��9K�9շ :b[:b[:׸ :��9n��9{�9���9L��9x   x   @��9Ok�9&}�9�N�9���9�9��9��9��9ʋ�9��9{M�9�~�9k�9���9���9���9���9�D�9��:��:C�:�0:�:ȳ:N�:�D�9?��9��9\��9x   x   ���99��9�C�9���9K�9��9{��9���90��9�I�9���9wD�9˶�9���9���9���9��93A :+:X�:i::�:N:�::�:L+:�@ :X��9?��9��9x   x   d�9�e�9@��9��9��9��9��9ζ�9���9l�9C��9�d�9��9��9mw�9|�9�E�9Z+:�*:Aw:��	:f
:��	:�v:*:�+:�E�9�{�9_z�9$��9x   x   ���9��9��9���9َ�9��9B�9]��99��9��9s��9���9���9v�9���99��9��:،:�w:R�
:�:Γ:��
:�w:e�:`�:���9���9M�9K��9x   x   *�9"�9��9;��9/�9m/�9 	�9w��9���9_#�9e��9��9���97`�9$��9��9��:(;:a�	:L�:O%:�:d�	:�;:��:C�9 ��9rc�9���98�9x   x   ��9|��9�Ľ9�H�9���9��9�F�9�ý9)��9s��9D|�9��9E�9�M�9�0�9?� :t�:�:�f
:E�:S�:�g
:�:D�:� :�1�97K�9�C�9���9�|�9x   x   ���9$f�9�޵9[!�9
>�9�"�9��9�g�9���9�>�9*$�9���9*B�9���9t��9�\:W2:t:��	:��
:��	:�:.2:f]:���9���9�C�9���9�$�9/=�9x   x   2��9V�9�N�9Kl�9Il�9�M�9(�99��9ٿ�9vD�9���9\>�9���9�Z�9W)�9]:��:�;:�w:�x:b<:��:�]:*�9�[�9V��9=�9h��9�E�9���9x   x   ���9�?�9�a�9�i�9fa�9�B�9��9 n�9Xk�9(��9m��9�i�9��9_[�9���9�� :X�:<�:+::�:��:j� :(��9�[�9�9�j�9(��9,��9Sj�96n�9x   x   d�9�F�9�M�9�N�9	D�9z�9ѱ�9��9��9�E�9Q��9�i�9���9J��9�/�9�9��:�,:-:3�:m�9�2�9k��9���9�j�9���9�D�97��9��9��9x   x   �:�9�V�9Q�9�X�9";�9��9J�9T5�9xI�94B�9���9=�9SC�9rN�9S��9��9�G�9�A :�G�9��9��9�K�9�C�95=�9%��9�D�9J�9�4�9�H�9��9x   x   d��92��9#��9G��9�\�9^Σ9!֪9�4�9���9���9k��9���9KC�9�a�9���9U~�9��9���9h}�9���9Sd�9/D�9��9\��9���9���9�4�9jת9Mϣ9�\�9x   x   �u�9G��9�w�9k5�9-��9�ϣ9HI�9��9�i�9�E�9�"�9h��9^��9F�9�{�9���9���9,��9�{�9B�98��9��9�$�9�E�9�i�9V�93H�9ϣ9���996�9x   x   ��9�9���9�5�9UZ�9z�9��9�m�9ľ�9�=�9d}�9��9���9��98��9���9Y��9���98��9ښ�9_�9d|�9�<�9R��9m�9Q��9�9\�9�5�97��9x   x   �!�9��9��9yl�9#�9�ͮ9]R�9�s�9���92�9�)�9�m�9��9*��9�9Y��9��9ם�9��9�m�9�(�92�9J��9r�9�S�9Ю9�9il�9���9��9x   x   s�9�:�9y�9Q��9@��9�l�93�9�9Ԯ�9V{�9m��9�*�9f|�9��9��9i�9\��9;~�9 ,�9ɾ�9�{�9��9���9��98i�9���9�9*�9y=�9��9x   x   9�9%�9Y�9��9^�9Ĵ9�9p�9#��9���9�g�9���9kj�9͎�9jQ�9ѐ�99j�9���93g�9��92��9,o�9��9�Ĵ9��9!�9�9`�9u��9b�9x   x   �k�9���9B�9�7�9�$�9/��9c��9>��9BL�9:��9D�9���9��9G��9*��9/��9���9�E�9��9�I�9,��9A��9f��9�$�9�4�9��9���9!l�9~J�9H�9x   x   ��9G��9��9�$�9��9��9�{�9W��9���9�i�9/+�9��9���9�a�9 ��9��9:*�9�h�90��9S��9�x�9O�9�9%�9I�99��9M�9���9��9ڎ�9x   x   ̮9Rk�9ô9���9n�9���9���9�#�9Vk�9�!�9��9�0�9�8�9:�9N1�9K�9#�9Uj�9"�9��9Y��9��96��9D´9(j�9�ή9��9��9@�9��9x   x   ~P�9��9��9���9{�9E��9���9�v�9���9���9q�9/j�9���9�g�9�9���9���9�w�9��9��9lz�9p��9J�9p�9�P�9}�9W�9O�9IT�9��9x   x   �q�9(��9�n�9$��9���90#�9{v�9}�95&�9�R�9��9#��9O��9���9�Q�9>%�9�|�9kw�9�"�9���9���9:m�9�9r�9���9 r�9�ո9�ָ9vr�9���9x   x   ���9ܬ�9���9
K�9���9�j�9;��9&�9�97��9tm�9	��9�j�9W��9<!�9O'�9���9�j�9���9K�9���92��9N��9~Q�9*=�9A��9iX�9���9C:�9vR�9x   x   0�9;y�9K��9��9�h�9/!�9G��9�R�9)��9�`�9��9���9�b�9��9yO�9S��9�"�9�g�9!��9���9*z�9�/�9�$�9�O�9���9��9��9���9_R�9�"�9x   x   '�9U��9f�9�B�9:*�9�9�9���9nm�9��9���9���9\k�9���9��96�9�)�9;D�9?g�9_��9�%�9��9Rf�9�9�9p�9!�9��9�7�9Ie�9��9x   x   k�9�(�99��9d��9��9j0�9�i�9��9��9���9���9H��9��9h�9�/�9w�9���9��9�(�9Al�9��9\�9`�9���9M��9-��9Ŭ�9�a�93�9���9x   x   ���9qz�9�h�9Ɍ�9 ��9�8�9���9e��9,k�9�b�9�k�96��9K��9�9�9���9���9k�9<{�9��9k��9��9��9(��9DU�9�}�9"T�9���9:�9d��9r��9x   x   ��9I��9v��9b��9ea�9�9�9�g�9A��9ƌ�9���9,��9uh�9,:�9O`�9���9��9
��9:��9��9���9���9�$�92=�9r��9$��9?=�9�%�9���9���9m��9x   x   D�9��9ZP�9���9���9g1�9^�9!R�9�!�98P�9t�9�0�9e��9���9�P�9�9R�9v�9�"�9`��9H�9�#�9iN�9���9�N�9y!�9H�9���9%%�9��9x   x   ���9I�9��9���9��9��9���9%&�9T(�9c��9C�9u�9���9���9^�9���9���9��9ќ�9��9��9��9���9���9o��9B��9)��9��9���9���9x   x   O�9���9�i�9���9�*�9�#�9���9�}�9���9�#�9*+�9���9,l�9��9��9��9���9��9���9~��9GU�9��9)��9��9aS�9΋�9���9���9���9���9x   x   ��9�}�9���9F�9yi�9bk�9(y�9�x�9\l�9�i�9�E�9���9�|�9���9��9���9d��9[��9���9*& :Dz:�):�*:{:Q& :)��9"��9���9���9��9x   x   ���9�+�9�g�9ў�9B��9e#�9���9�$�9���9+��9Gi�9�*�9��9���9($�9��9m��9���9n� :}:��:^ :Ŝ:}:>� :��9���9W��9)&�9`��9x   x   �m�9��9���9�J�9���9���9���9���9RM�9?��9���9�n�9���9���98��9���9���9�& :<}::��:��::6}:f& :��9���9
��9���9���9x   x   >)�9&|�9!��9w��9oz�9M��9�|�9��9@��9�|�9�(�9���9���9��9DJ�9���9�V�9�z:�:��:j:��:�:M{:1W�9۩�9.J�9z��9%��9��9x   x   �2�9���9]p�9ɑ�91�9�9ِ�9�o�9���9�2�9��9T�9��9�'�9&�9S��9��9E*:� :��:��:b:+: �9��9�&�9�%�9��9S�9&��9x   x   ���9���9	�9��9�9���9��9���9N��9�'�9�i�9<c�9P��99@�97Q�9:��9`��9�+:|�:�::�:@+:1��9:��9�N�9tA�9���9%e�9�h�9,%�9x   x   �r�9��9/ƴ9�&�9F'�9�Ĵ9+�9�t�9�T�97S�95=�9��9�X�9���9���9m��9b�9%|:�}:�}:�{:x�9d��9%��98��9�W�9���9^;�9bU�9YU�9x   x   �T�9tj�9I�9�6�9|�9�l�9�S�9���9d@�9���9�!�9���9A��9y��9�Q�9F��9�U�9`' :� :' :'X�9���9#O�9W��9K��91��9�#�9���9$?�9���9x   x   �Ю9杫9��9��9o��94Ѯ9��9*u�9���9}��9��9���9�W�9�@�9�$�9��9L��9I��9���9g��9̪�9�'�9�A�9X�90��9t�9g��9��9w�9΀�9x   x   ��9��9��9F��9l�9��9�Y�9ظ9�[�9D��9T#�9?��9
��9�(�9
K�9���9���9,��9:��9���9K�9l&�98��9���9�#�9U��9*]�9ٸ9�W�9��9x   x   m�9+�9��9�m�9���9��9��9dٸ9���9/��9;�9�d�9��9���9���9}��9Â�9���9˞�9��9*��9��9Ae�9T;�9���9��9�ظ9]�9��9���9x   x   S �9E>�9� �9�K�9l�9Y�9�V�9u�9&=�9dU�9Yh�9M�9q��9���9�'�9���9���9���9R'�9���9���9u�9�h�9 U�9�>�9�v�99W�9z�97�9�K�9x   x   ��9i�9c�9=I�9m��9��9��9���9U�9f%�9Ͻ�9P��9+��9��9� �9���9���9��98��9c��9��9��9�$�9�T�9c��9,��9�9T��9�K�9�c�9x   x   �J�9��9$��9�}�9C_�9�9x�9�U�9Oi�9�l�9'�98�9��9���9���9�v�9���9���9���9�9�9�%�9�k�9Oj�98T�9bz�9@�9�^�9�}�9��9��9x   x   ��9��9<$�9�^�9�l�9�6�99��9~3�9���9ds�9��9j�9���9��9%D�9
D�9��9~��96�9��9\t�9���9<4�9z��95�9$m�9�^�9V$�9���9p�9x   x   ���9�#�9%��9h�9�1�9
�9��9j�9Ͱ�9���9<)�9T��9թ�9�l�9O��9Rm�9���9���9L)�94��9i��9h�9��9��9�2�9��9��9�#�9ؠ�9\�9x   x   �|�9k^�9 �9Ȉ�9I��9�/�9���9���9 ��9=��9��9���9���9���9���9���9���9T��9k��9���9l��9��9O.�9L��9n��9L�9M^�9�|�9]��9���9x   x   :^�9-l�9i1�9��9t��9���90�9���9��9�W�9�p�9!��9�7�9���98�9��9�p�9�V�9ɭ�9���9�-�9���9W��9���9\2�9�k�9�^�9��96��9�9x   x   ��9�5�9D�9X/�9A��9Ԛ�9ew�9+F�9t��9���9�1�9@��9 ��9δ�9&��9�1�9���9���9�D�9�w�9���9���9�-�9�9�4�9��9���9�Ѳ9�Ҳ9���9x   x   �v�9센9��9���9�/�9,w�9��9���9��9��9!��9s��9P�9T��9u��9!�9p��9&��9n��9�v�9�-�95��9x�9C��9�w�9	�95��9���9���9��9x   x   T�9�1�9�h�9���9��9�E�9���9�c�9���9	?�9�v�9W�9_�9�w�9�>�9���9Vb�9���9�D�9���9���9�g�941�9;S�9�߾9۽94\�9<]�9�۽9߾9x   x   mg�9	��9}��9��9`��9���9���9{��9�9�.�9��9W&�9���9�-�9(�9��9���9���9Q��9ޝ�9s��9I��9�h�9_+�9gF�9��9��9���9�D�9�,�9x   x   �j�9�q�9L��9��9�V�9S��9k�9�>�9�.�9*��9�A�9�A�9���9�.�9N=�9�9U��9LW�9���9:��9�r�9�h�9��9���9�|�9�I�9'I�9B~�9���9~��9x   x   %�9R��9�'�9��9�o�91�9���9�v�9���9�A�9�V�9aA�9���9�w�9e��90�9�o�9y��9d)�9ʌ�9�%�9<��9���9cj�9iF�9�C�9WF�9�h�91��9���9x   x   6�9��9���9���9i��9���9/��9?�9d&�9�A�9sA�9	'�9��9G��9���95��9���9���9	�9H6�9ҏ�9;��9��9�C�9�a�9Eb�9XD�9��9U��9΍�9x   x   &��9���9���9���9E7�9ȳ�9 P�9m�9"��9���9���9
�9�P�9���9�5�92��9��9���9@��9���9js�9�C�9w��9qK�9�s�9JJ�9T��9_A�9�s�9���9x   x   ���9.�9�k�9���9���9���9a��9�w�9!.�9
/�9x�9���9ȴ�9<��9���9_j�9��9l��9c~�9]#�94��9��9Ƴ�9�#�9�$�9g��9G��9���9� �9}�9x   x   ��9�B�9v��9Q��9�7�90��9���9k?�9��9�=�9���9Y��9!6�9��91��9ZC�9���9�>�9֯�9i��9u��9M�9t4�9���9�3�9�K�9o��9S��9z��9�?�9x   x   \u�9C�9�l�9���9&��9 2�9��9���9ވ�9��9�0�9���9���9�j�9�C�9Dr�9��9V��9U��9���9s��9!G�9��9��9�H�9���9D��9U��9���9��9x   x   ���9	�9m��9���9-q�9m��9?��9Jc�9���9v��9�p�9���9ݫ�9n�9X��9e��9���9�}�9v��9���9a�9E��9V��9��9,�9���9���9=~�9Y��9��9x   x   ��9$��9|��9���9JW�9���91��9���9��9�X�9���9���9ʏ�9z��9�?�9���9*~�9n��9�x�9j��9��9���9G��9���9U��9�x�9���9�~�9���9�?�9x   x   1��9,�9�)�9���9���9�E�9���92F�9��9���9+�9��9Ą�9��9��9>��9��9Iy�9lR�9!7�9��9a��91�9�7�9R�9z�9���9^��9`��9�~�9x   x   �9�9A��9���9Z��9��9�x�9Kx�9���9���9*��9Ď�948�9a��9	%�9���9ɚ�9���9��9q7�9���9�'�9�)�9��9%7�9M��9��9;��9n��9�#�9���9x   x   �%�9�t�9/��9���9-/�9:��9{/�9���9���9�t�9�'�9���9�u�9"��9>��9��9��9��9c	�9(�9���9!(�9�	�95��9��99��9���9a��9�u�9m��9x   x   \l�9���9i�9?��9`��9���90 �9�i�9���9�j�9���9���9F�9L��9O�9�H�9̄�9.��9S��9*�9b(�9N��9ܼ�9L��9GJ�9�O�9��9�E�9Q��9)��9x   x   �j�95�9��9�/�9���9�/�9��9�3�9.k�9z��9U��9+�9��9<��9�6�9��9�9���9K�9���9d
�9��9<�9;�9%5�9��9���9h�9���9=��9x   x   �T�9d��9'�9Ϊ�9^��9�9|��9�U�9�-�9y��9-m�9�F�9#N�9&�9��9��9߄�9��99�98�9ס�9���9g�9���9�&�9�M�9wF�9|l�9s��9�/�9x   x   {�9�5�94�9���9.4�9�6�9z�9i�9I�9��9?I�9yd�9Rv�9�'�9V6�9�J�9)�9��9fS�9_��9J �9�J�9d5�9�&�9�u�9e�9I�9V��9�G�9��9x   x   �9n�9��9��9�m�9��9S�9�ݽ9���9�L�9�F�9*e�9M�9��9#N�9B��9���96z�9a{�9��9���9P�9*��9N�9e�9yF�9�L�92��9#޽9��9x   x   �_�9�_�9W��9�_�9C`�9���9s��9�^�9���9�K�9,I�9+G�9��9���9���9���9���9���9��97��9A��9q��9���9�F�9
I�9�L�9b��9�_�9* �9䗳9x   x   U~�9-%�9�$�9/~�9��9�Ӳ9���9�_�98��9��9gk�9��9�C�91��9���9c��9��9��9���9A��9��9�E�9��9dl�93��9��9�_�9ª�9tղ9�9x   x   ���9���9ġ�9���9���9�Բ9���9޽9/G�9S��9���9���9Tv�9�"�9���9`��9��9���9U��9{$�9�u�9n��9���9:��9�G�9�ݽ9���9Eղ9+��9�9x   x   ��9��9�9��9b�9.��9��9�9�.�9���9��9��9/��9�9\A�9���9X��9�@�9A�9��9���9��9��9%/�9o�9E�9n��9��9Ҋ�9��9x   x   p��9I1�9���9�	�9i8�9��9���92`�9ga�9�T�9��9�.�9>��9�H�9���9\y�9��9[I�9��9[0�9+�9�T�9�`�9_�9��90�99�9�	�9^��9[1�9x   x   1�9!�9��9���9��9��9E�9���9���9�-�9q]�9J��9���9B��9���9���9��9���9���9�\�9�.�9���9���9C�9*�9��9^��95�9m �9�0�9x   x   >��9^�9��9Ӷ9�@�9�"�9_\�9���9d
�9� �9���9d��9�9a��9��9Ս�9#�9Q��9���9Y!�9r	�9ú�9*^�9�#�9�@�9�Ҷ9_�9��9 ��9G6�9x   x   ��9;��9�Ҷ9��9
�9G��9���9u��9���9�0�9�C�9Ͻ�9nl�9]P�9P�9?m�9Ż�9�C�9F0�9=��9ɿ�9��9���9	�9,��9�Ҷ9
��9z�9�>�9�>�9x   x   �7�9M�9�@�9�	�9a<�9'��9vU�9s��9�A�9�G�9d��9	��9.��9iI�9��9*��9��9G�9C�9���9�T�9a��9!>�9�	�9<?�9��9�8�9)�9�д9�)�9x   x   r�9�9="�9���9��9���9��9 "�9���9�f�9�W�9ް�9vl�9�l�9+��9sW�9�e�9��9a!�9��9���9���9���9�"�9�9X�9�9�O�9�N�9��9x   x   d��9�C�9�[�9���9U�9��9Z��9�=�9b��9�j�9 ��9T��9
�9ܾ�9���9�i�9��9+=�9���9Q�9�T�9���9�[�9oD�9��9AI�9���9�D�9���9eH�9x   x   �^�9���9���9���9���9�!�9�=�9�;�9���9�]�9+[�9Y��9���9Z�9�^�9?��9W:�9u=�9� �9���9���9ɻ�9M��9�]�9�3�9�h�9O��9���9�i�9S3�9x   x   �_�9T��9I	�9��9A�9&��9��9���9�,�9o�9֬�9���9h��9��9f,�9���9��9k��9�B�9B��9I�9L��9�a�9Na�9��939�9L�9�7�9���9�a�9x   x   BS�9�,�9��90�9G�9f�9�j�9�]�9e�9��9$��9���9p��9��9�]�9�i�9<e�9tG�9�-�9� �9u,�9,Q�9{��9�9���9���9ڒ�9��9T�9���9x   x   ) �9\�9���9C�9���9W�9���9[�9ͬ�9'��9&��9��94��90[�9>��9�V�9���9�C�9���9[�9��9ٰ�9���9�[�9�Q�9Q�9�O�9�[�9���9���9x   x   �,�9���9A��9��9k��9s��9$��9N��9���9���9,��9��9&��9L��9��9���9��9q��9���9X,�9d�9<��9
��9��9t�9��9���9���9Ѡ�9Od�9x   x   ���9���9�9�k�9���9$l�9��9���9���9���9Y��9:��9��91l�9���9�l�9E�9���9S��9�y�9�7�9{��9#k�9���9N��9��9�i�90��9�7�9{�9x   x   9G�9��9w��9�O�9
I�9�l�9��9;Z�9��9P�9w[�9���9Vl�9�I�9�O�9V��9-��9�E�9���9l�9^B�9m<�9���95N�9�N�9E��9�<�9mB�9�9I��9x   x   Z��9���9�
�9�O�9���9/��9��94_�9�,�9O^�9���9Y��9���9�O�9N�9���9���9���9���9t��9xO�9q�9�,�9\u�9�+�9�q�9N�9��9e��9��9x   x   Qx�9���9I��9�l�9*��9�W�9�i�9���9j��9|j�9�W�9E��9um�9���9���9�u�9�9���9�+�9#R�9��9PE�9N��9���9�D�9��9�Q�9�+�9ۼ�9��9x   x   O��9���9��9Ż�9U��9af�9���9;�9���9"f�9y��9Ż�9�9���9J��9C�9�S�9�o�9�8�9U��9b�9�}�9��9c�9�`�9���9�7�9Gp�9�S�9b�9x   x   �H�9h��9H��9D�9�G�9(��9>�9w>�9~��9�H�9�D�9���9~��9�F�9���9x��9&p�9u��9R��9�O�9s�9���9��9q�9�O�9x��9���9=p�9���9���9x   x   ���9���9���9�0�9�C�9C"�9��9�!�9�C�9/�9!��9��9���9���9���9i,�99�9���9���9�C�9*��9�8�9
��9'D�9���9���9�8�9f+�9���9x��9x   x   F0�9�\�9�!�9��9���9��9��9k��9̞�9q"�9�\�9�-�9T{�9��9���9&S�9��9/P�9�C�9	^�9�p�9�q�9P[�9�C�9�P�9���9pT�9D��9�9M{�9x   x   L�9�.�9
�9���9�U�9��9?V�9O��9
�9<.�9��9�e�9�9�9�C�9�P�9�9	c�98�9���9#q�9�9^q�9��9��9c�9��9�O�9:C�9�9�9�e�9x   x   �T�9%��9���9��9���9t��9r��9���9/��9$S�9ܲ�93��9f��9?>�9�r�9�F�9�9���9�9�9r�9�q�9H9�9���9n�9?G�9�r�9v?�9��9��9m��9x   x   Za�9���9_�9��9�?�91��9�]�90��9�c�9���9ʅ�9.��99m�9{��9�.�9���9m��9F��9��9�[�9���9���9���9���9�.�9c��9�k�9���9���9t��9x   x   �_�9�C�9�$�9I
�9d�9~$�9@F�9�_�9uc�9D�9^�9L �9ü�9TP�9Ww�9v��9��9��91E�9�D�9C�9��9���9�x�9P�9@��9��9�^�9��9�d�9x   x   ���9��9�A�9g��9�@�9��9���9�5�9D��9���9�S�9��9���9Q�9�-�9�F�9�b�9�P�9��9eQ�9�c�9�G�9�.�9P�9���9N�9R�9���9���9�6�9x   x   ��9��9�Ӷ9�Ӷ9B�9�9(K�9k�9`;�9��9tS�9��99��9n��9�s�9��9���9���9���9q��9p�9(s�9���9R��9O�9�T�9/��9�<�9�i�9I�9x   x   �9�9��9X�9>��9):�9��9q��9X��9p�9��9R�9�9�k�9"?�9�O�9�S�9T9�9��9�9�98U�9hP�9�?�9�k�9��9R�9"��9��9���9���9��9x   x   K
�9��9��9�	�9`*�9KQ�9<F�9���9�9�9/��9^�9!��9S��9�D�9���9V-�9�q�9hq�9O,�9��9�C�9R��9���9�^�9���9�<�9���9+C�9�P�9`*�9x   x   ���9� �9ﭰ9�?�9=Ҵ94P�9-��9Zk�9���9\�9��9��9�9�9 �9��9f��9�T�9���9Y��9��9�9�9,��9���9��9G��9Qi�9x��9�P�9�Ҵ9�?�9x   x   �1�9�0�9�6�9�?�9�*�9�9�I�9�4�9�c�9���9���9)f�9�|�9���9���9��9u�9l��9���9�{�9�e�9J��98��9md�9o6�9�H�9��9*�9a?�9�6�9x   x   �Ǵ9R.�9�b�9�R�9���9�7�9.��9���9���95��9��9�9�9�97�9b��9���9���9j8�9Q�9l:�9���9���9:��9���95��936�91��9�R�9�e�9�.�9x   x    .�93�9�u�9J��9r`�9f��9�E�9J�9'��9k��9�9v�9Yg�9W�9���9j��9�9f�9��97�9Ҧ�9P��9E�9pD�9q��9`�9u��9Jt�9 �9�.�9x   x   Qb�9yu�9�)�9�w�97L�9�|�9���95��9��9ml�9�a�9���9��9��9BN�90��9���9���9_b�9�k�9�9��9K��9�}�9GK�9�v�9�+�9av�9�c�9d�9x   x   :R�9�9gw�9Ͻ9��9��9���9�4�9�`�9�G�9l��9���9�2�9+��9���9�3�9���9K��9�G�9�`�9d5�9���9���9:��9ҽ9;v�9���9�R�9ư�9���9x   x   ��9�_�9�K�9��9�=�9��9�9��9y��9�)�9�,�9��9!��9j��9���9(��9,.�9�)�9د�9���9��9��9N?�9���9�I�9zb�9���9��9�ӹ9X�9x   x   7�9���9<|�9©�9��9���964�9��9��9��9��9���9zF�9>F�9O��9��99�9I�9ܰ�9�4�9��9,�9��9�|�9���9�4�9�7�997��9�8�9x   x   ��9�D�9���9#��9��94�91]�9w�9�L�9-��9%�9
��9z��9~��9A�9���9�N�9v�9
]�9�3�9
�9B��9J��9$E�9���9F��9.0�9���9�1�9���9x   x   ���9C�9g��9^4�9���9گ�9�v�9>�9�p�9ӏ�9�L�9���9o��9K�9ڐ�9q�9f�9�w�9��9���9�2�9��9��9D��9W��9�,�9���9V��9�-�9���9x   x   ���9
��9 �9`�9��9^�9�L�9�p�9�q�9-�9�9���9M��9�,�9fq�9_p�9�M�9[�9K��9{`�9��9[��9?��9��9W|�9� �9?�97�9�}�9��9x   x   ���9>��9vk�9
G�9@)�9��9���9���9-�9!��9D��9n��9���9-�9���9��9��9f)�9�E�9�k�9���92��9~l�9���9��9��9ȏ�9��9���9em�9x   x   ���9��9�`�9���9�+�9���9��9�L�9���9L��9��9]��9z��9LL�9��9��9D-�9o��9a�9�9	��9��93j�9L�9bG�9�.�9�D�9N�9,k�9��9x   x   ,8�9L�9���9��9���9H��9ؽ�9���9���9{��9m��9���9V��9پ�9���9E��9���9��9_�9_8�9d�9Y��9@��9���9���9���9���9e��9���92g�9x   x   ��9Jf�94��9Y2�9���9?F�9Y��9w��9m��9י�9���9n��9��9�E�9���9�3�9;��9�e�9]�9]��9�V�9��9�F�9Έ�9���9ۈ�9�E�9���9zT�9���9x   x   �5�9`
�9R��9���9��9#F�9~��93K�9�,�9L-�9�L�9��9�E�9t��9���9H��9�
�97�9S�97s�9p�92�9���9��9��9z��9�0�9o�9<u�9cU�9x   x   Y��9���9�M�98��9g��9T��9j�9��9�q�9���9^�9���91��9��9mN�9���9$��9�0�9��9�E�9s|�9bq�9�9�,�9{�9�s�9g{�9�G�9���90�9x   x   ���9���9���9�3�9%��9��9"��9�q�9�p�9���9���9Ⱥ�9W4�9���9���9���9b"�9�@�9	=�9���9�Z�9]�9���9���9/Z�9^[�9���9�<�9�C�9�!�9x   x   S��9�
�9`��9���9Y.�9��9O�9��9FN�9_�9 .�9���9ҿ�9�9���9�"�9(��9�8�9}��9�f�9���9��9t�9��9���9�f�9��99�9���9�"�9x   x   �7�9�e�9���9y��9 *�9��9�v�9�x�9>�9N*�9[��9���9Zf�9�7�961�9NA�99�9k�9or�9_�9|��9gv�9er�9i��9�^�9�r�9x�9�8�9@D�9�0�9x   x   �9��9�b�9=H�9e��9���9�]�9��9f��9�F�97b�9y�9`�9T�9���9�=�9��9�r�9���9N��9+��9�X�9���9���9���9gr�9���9�<�9���9T�9x   x   ^:�9\�9Fl�9ta�9���9�5�9�4�9���9�a�9@m�9d�9�9�9���9Qt�9�F�9x��9�g�9{_�9���9�v�9�K�9HK�9�s�9���9�_�9
g�9,��9}H�9�w�9���9x   x   ���9��9�96�9�	�9���9J�9P4�9�9��9���9�e�9WX�9pq�9�}�9�[�9R��9��9���9�K�9���95L�9f��9"��9���9�\�9n}�9�n�9�V�9g�9x   x   ���9���9�9{��9��9T�9���9k��9���9���9���9��9���9�3�9�r�96^�9��90w�9Y�9�K�9ZL�9X�9�t�9��96]�9!r�9@5�9���9��9G��9x   x   ���9��9��9f��9h@�9Z��9���9��9���9:n�9�k�9���9VH�9f��9��9��9��9Ss�9E��9t�9���9�t�9��9���9a	�9���9�F�9���9'k�9pp�9x   x   Z��9E�9Q~�9E��9Г�9~�9�F�9���9_�9���9�M�9���9���9��9f.�9��9Q��9v��9i��9|��9���9U��9���9�.�9��9ċ�9`��9kP�9���9��9x   x   ���9 ��9%L�9ӽ9�J�9���9���9 ��9#~�9Ļ�9HI�9���9t��9s�9�9�[�9B��9�_�9���9C`�9f��9�]�9�	�9��9[��9z��9�F�9x��9 ~�9:��9x   x   �6�9�`�9�w�9Aw�9�c�9>6�9���9:.�9�"�9���9h0�9���9���9@��97u�9�\�9h�9�s�9Is�9�g�9]�9nr�9���9ڋ�9u��93�9d��9�$�9H,�9 ��9x   x   ���9 ��9�,�9���9(��9=9�9�1�9B��9 
�9���9�F�9��9�G�9�2�9 }�9,��9H��9��9a��9���9�}�9�5�9�F�9p��9�F�9Q��9��9���984�9�9�9x   x   S�9�t�9w�9oS�9��9<��9:��9���9� �9ʺ�9�O�9.��9���9�p�9I�9>�9F:�9�9�9�=�9I�9�n�9��9���9dP�9d��9�$�9���9}��9���9��9x   x   f�9w�9-d�9���9�Թ9j��9M3�91/�9&�9;��9�l�9Z��9V�9�v�9���9E�9���9E�9Q��9�w�9!W�90��9k�9���9�}�9,�9	4�9x��9ع9걷9x   x   �.�9/�9��9[��97�9:�9��9+��9X�9�n�9���9�h�9)��9�V�9T1�9#�9�#�9�1�9�T�9Ȳ�9g�93��94p�9V�9���9���9�9�9��9ȱ�9>�9x   x   ��9�
�9��9��9�Ծ9�w�9�u�9���9��9g�9o��9cR�9y��9Lc�9O{�9Q��9�x�9+e�9���9VR�9)��9�g�9�9��9s�9�t�9�׾9��9d�9�
�9x   x   �
�9#��9A�9���9���9
��9���9���9���9/��9���9�-�9��9�q�9 �9"�9r�9�9�,�9y��9:��94��9���9��9:��9���9ܲ�9J߻9㥺9�9x   x   p�9�9�K�9�5�9;��9�)�9x�9���9y��9���9"�9l�9k��9��9��9���9���9R�9��9ԕ�9��9���9��9*�9\��95�9�O�9)�9��9C��9x   x   ���9C��9�5�9�"�92s�96��9���9�K�9%��9X@�9]R�9���9K�9���9���9��9)��96Q�9�@�9Z��9�J�9���9"��9�q�9&�9�3�9ⰽ9橼9��9��9x   x   �Ӿ9��9��9s�9ɝ�9]��9�T�9h��9$��9���9���9��9e��9���9���9���9P��9���9���9B��9�U�9���9���9�r�9ˉ�9��9�Ծ9B�9�ܽ9��9x   x   �v�9r��9�)�9���9A��95�91#�91�9�
�9���9���9x��9#Q�9SP�92��9���9��9k	�9�2�9�#�9g�9���9=��9�)�9q��9@u�9��9�7�96�9-��9x   x   �t�9���9��9N��9[T�9#�9���9���9��9�V�9�D�9���9	�9K��9HE�9�U�9��9ƒ�9p��9t"�9pV�9��9��9.��9[r�9M��9��9���9��9��9x   x   ǹ�9ѽ�9 ��9>K�9��9�0�9���9���9� �9.��9|��9���9���9Q��9���9
 �9���9|��92�9���9�I�9���9"��9���93��9Ff�9- �9B�9h�9��9x   x   ��9��9���9���9���9I
�9X�9� �9���9o]�9V��9��9���9�]�9x��9���9��9	�9n��9��9��9\��9k�9s�9 ��9B��9���9���9
��90r�9x   x   �e�9A��9��9�?�9��9_��9V�9��9i]�9°�9��99��9M��93\�9:��9�V�9ʫ�9���9�?�9̕�9��9�g�9���9���9�\�9�?�9C�9n[�9k��9I��9x   x   N��9���9V�9�Q�9/��9���9�D�9b��9L��9��9���97��9(��9���9_C�9x��9o��9�P�9�9���9���9�\�9&8�9�!�9�9y�9��9�$�9�9�9h[�9x   x   KQ�9�,�9��9U��9���92��9���9���9���9=��9A��9��9���9r��9��9���9E��9!�9k,�9R�9W}�9��9���9���9q��9���9j��9[��9Þ�9/��9x   x   n��9��9���9��9��9�P�9�
�9���9���9d��9=��9���9�	�9^P�9X��9&�9���9�9X��99�9Ѳ�9��9�t�9֧�9v��9T��9�u�9�$�9l��946�9x   x   Yb�9�p�9���9<��9���9;P�9J��9k��9�]�9o\�9���9���9wP�9Z��9��9؆�9r�9�d�9$\�9�8�9��9 ��9	�9�V�9�U�9��9ש�9�9y<�9�^�9x   x   xz�9b�9���9<��9���91��9iE�9���9���9���9�C�9Y��9���9,��9���9��9�v�9@��9e*�9�L�9�M�9��9ƌ�9&��9���9�9�M�9:N�9�%�94��9x   x   ���9y!�96��9��9���9���9V�9f �9W �9(W�9���9��9��9��9 �9���9R��9]M�9$��9AS�9�s�9n;�9P��9t��9�7�9�s�9�R�9_��9R�98��9x   x   �w�9�q�9]��9��9v��9;��9��9���9a�9l��9��9���93��9r�99w�9��9��9���9���9�9�B�9.��9Q=�9p��9D�9��9��9Y��9���9���9x   x   �d�9��9J�9VQ�9���9�	�9T��9"��9�	�9N��9�Q�9��9��9he�9���9�M�9���9��9���9��9���9l,�9)�9��9N��9��9X�9&��9�P�9s��9x   x   p��9�,�9�95A�9j��9D3�9!��9�2�9F��9�@�9��9J-�9-��9�\�9
+�9���9	��9%��9r��9�n�9R[�9H��9I^�9o�9M��9D��9���9���9�&�9-]�9x   x   LR�9���9��9���9޸�9�$�9P#�9u��9��9ܖ�9���9!S�9 :�9�9�9dM�9�S�9��9<��9�n�9i��9�z�9�y�9N��9�n�9i��9P�9�Q�9O�9�>�9<7�9x   x   <��9}��9|��9�K�9pV�9@�9fW�9�J�92��9H��9��9�~�9���9��9�N�9�t�9�C�9��9�[�9�z�9t��9R{�9N^�9���9�C�9v�9!P�9��9���9��9x   x   �g�9���9 ��9���9}��9���9��9���9���9�h�9^�9U��9>!�9O��9��9`<�9���9-�9���9Oz�9v{�9��9�+�9���9P:�9?�9Ȯ�9$�9���9(\�9x   x   Z�9��9M�9���9���9R��9�9h��9��9��9�9�94��9"v�9[�9���9f��9A>�9�)�9�^�9���9�^�9�+�9x>�9{��9L��9�9u�9���98�9��9x   x   H��9���9�*�9�r�9vs�9�*�9r��9���9ut�9/��9/#�95��9G��9�W�9r��9���9j��9��9�o�9<o�9	��9���9���9���9�V�9��9��9�&�9���9r�9x   x   {s�9Ħ�9��9�&�9Њ�9���9�s�9���9���9^�9��9���9���9W�9���9�8�9$E�90��9��9���9SD�9�:�9q��9�V�9��9���9��9|\�9���9���9x   x   9u�9L��9�5�9�4�9��9\v�9���9�g�9���9A�9
�99��9թ�9�9n�9$u�9��9���9 ��9��9qv�9~�99�9���9���9>�9�A�9ϣ�9Uf�9��9x   x   �׾9c��9^P�9���9�վ96��9�9�!�9#��9�D�9a�9���91w�9B��9KO�9�S�9��90�9M��9+R�9P�9���9u�9!��9��9�A�9Տ�9� �9��9���9x   x   W��9�߻9��9���9,�9�8�9��9� �9��9�\�9$&�9���9!&�9l�9zO�9z��9Q��9���9e��9�O�9�9H$�9���9s&�9o\�9���9� �9O��9�6�9*�9x   x   ��9E��9 �9��9�ݽ9�6�9��9Hi�9X��9ŝ�9�:�9#��9���9�=�9�&�9S�9���9�Q�9.'�9?�9���9��9 8�9���9o��9-f�9��9�6�9��9*�9x   x   �9_�9���9��9c�9��9��9-��9`s�9���9�\�9j��9e7�9�_�99��9��9B��9��9�]�9q7�9���9\�9���9�q�9R��9���9:��9��9�9T��9x   x   2��9��9�ž9�9-��9A�9���9�8�9J��96��9G�9���9~o�9��9z��9w�9z��9���9op�9}��9�F�9��9\��9�:�9���9v�9��9W�9Ⱦ9��9x   x   ��9c�9��9���9B��93�9��9�	�9���9�#�9�m�9�f�9���9��9��9���9��9B��9pf�9Hn�9%$�9���9�	�9��9u�9d��9���9�~�9�}�9���9x   x   �ž9��9���91;�9s�9�J�9���9�9vg�9٥�9,��9H�9݌�9}T�9���9�S�9���93I�9��9g��9/g�9r�9Z��9�I�9��9�:�9���9���9�ž9J��9x   x   ��9���9;�97��9*��9���9���9��9�@�9�1�9���9�1�9��9��9.��9W�9,2�9���9�1�9ZA�9��9��9J��9Z��9���9:�9E��9��9���9���9x   x   ���9���96�9
��9j�9_�9�U�9�E�9"�9n��9�$�9m+�9���9���9���9C*�9�$�9���9�!�9rE�9�V�9�]�9*i�9���9�9���9���9.O�9[�9zO�9x   x   ��9��9J�9[��9�^�9��9S��9Rt�9���9�N�93\�9e�9�}�9~|�9�9u]�9�M�9��9�u�9���9��9�_�9���9�J�9,�9	�9h�9��9J�9�i�9x   x   ٓ�9n��9'��92��9�U�9:��9�;�9���9���9���9���9�9�<�9��9}��9z��9d��9��9�;�9{��9�T�9-��9d��9���9}��9���9�m�9I�9�n�99��9x   x   8�9��9��9|�9�E�9"t�9���9���9Ց�9�H�9���9��9}�9���9I�9i��9m��9A��9�u�9�F�9��9�9f�9*9�9���9�#�9���9���9�$�9ʍ�9x   x   h��9Р�9�f�9D@�9("�9���9���9ˑ�9�1�9���9{��9;�9i��9\��9�1�9	��9Q��9{��9 �9q@�9+f�9֡�9���9~n�9�9���9Q��9���97�9�n�9x   x   M��9 #�99��91�9��9�N�9���9�H�9���9���9x�9��9-��9I��9�J�9���9�M�9���9�1�9ͥ�9"�9N��9�R�9�	�9{��9��9���9��9��9�R�9x   x   "F�9 m�9���9Y��9C$�9�[�9ِ�9���9s��9|�9o$�9��9B��9���9D��9$]�9#�9��9v��9�m�9<F�9/�9��9���9���9���9��91��9��9�9x   x   ӈ�9�e�9iG�9r1�9+�9 �9��9��94�9��9��9B
�9��9��9 �9+�9�1�9I�9>e�9ǈ�9`��9<��9��9I��9�9��9{��9���9���9���9x   x   �n�9%��9L��9|�9V��9o}�9�<�9|�9w��9D��9R��9��9�;�9�|�9q��9��9?��9���9�n�9���9+E�9���9���9!�9u�9p�9���9ԟ�9ID�9+��9x   x   X��9K�9�S�9���9���9f|�9��9���9{��9r��9���9��9�|�9n��9���9T�9��95��9���9�R�9/��9G�9���9�97�9���9�}�9B��9$T�9P��9x   x   Ѻ�9f��9,��9��9���9�9���9LI�9�1�9�J�9���9\�9���9Γ�9u��9Ǟ�9k��9���9@��9���9���9�F�9���9H��9E��98H�9���9h��9���9���9x   x   �
�9D��9�S�91�9H*�9�]�9���9���9[��9���9~]�9o+�9
�9QT�9ߞ�9��9�y�9���9�+�9�N�97�9=��9)�9(�9���9�6�9�M�9+�9���9xx�9x   x   
��9D�9���9$2�9%�9�M�9���9ݦ�9���9qN�9�#�9b2�9���9 �9���9z�9m/�9���9JH�9ۈ�9z�9�
�9�;�9�9N{�9	��9�I�9)��9S.�9]{�9x   x   z��9��95I�9���9��9j��9~��9Д�9��9#��9���9J�9!��9���9Q��9���9��9s��9V<�9'��9�a�9G��9N��9/`�9m�9�;�9���9���9���9`��9x   x   Ep�9Zf�9��952�9�!�9\v�9<�9?v�9� �9U2�90��9�e�9[o�9H��9���9;,�9�H�9{<�9h��9��9k��9I�9���9C�9���9';�9J�91-�9j��9ӝ�9x   x   r��9]n�9���9�A�9�E�9)��9.��9�G�9FA�9���9�n�9���9���9bS�9h��9iO�9>��9o��9��9p$�9n��9���9�"�9��9Y��9_��9�L�9M��9�V�9���9x   x   �F�9W$�9�g�9J�9UW�9��9sU�9l�9g�9#�9<G�9V��9F�9 �9n��9�7�9�z�9	b�9���9���9r��9ܮ�9s��9�`�99z�9�9�92��9���9E�9��9x   x   ��9��9��9���9u^�9�`�9��9	�9��9`��9G�9L��9��9D��9�G�9
��9��9���9��9ݭ�9���9N
�93��9��9��9�E�9���9P��9|��9�9x   x   ���91
�9ܢ�9��9�i�9���9]��9v	�9���9�S�9�91��9���9���9���9�)�9<�9���9��9<#�9���9I��9{;�9[)�9���9���9���9���9��9�U�9x   x   !;�9i��9xJ�9 ��9q��9�K�9���9@:�9�o�9�
�94��9~��9T�9&�9P��9)�9��9�`�9��9�9�`�9��9m)�9���9�9��9���9Q��9�	�9!n�9x   x   ���9��9m�9���9��9(�9���9Ԏ�9I�9���9��9S�9��9[�9W��9���9-|�9!��9+��9Ɓ�9�z�9Q��9��9�9$�9b�9���9���9
�9��9x   x   ��9���9S;�9�:�9a��9��9���9�$�9���9X��90��9��9��9���9II�9�7�9��9�<�9�;�9݉�9�9�9�E�9���9��9_�9v��9���9���9�#�9L��9x   x   c��9Q��99��9���9���9i�9�n�9	��9���9���9D��9���9���9�9���9�N�9qJ�9G��9�J�9M�9}��9�9���9���9���9���9-��9���98o�9�i�9x   x   ��9�~�9��9k�9�O�9��9�I�9���9��9=��9c��9��9 ��9^��9l��9�+�9���9%��9�-�9���9���9p��9���9A��9���9z��9���9K�96�9�O�9x   x   UȾ9~�9ƾ9��9�9�9no�9�%�9K	�9��9��9���9dE�9&U�9���9���9/�9F��9���9W�9*E�9���9��9�	�9�	�9�#�9o�9-�9��9��9x   x   ,��9��9���9��9P�9Aj�9
��9���9�o�9�S�9�9���9&��95��9���92y�9�{�9���9��9���9/��9��9�U�9�m�9ӎ�9��9�i�9mO�9먿9t��9x   x   ���9��9g��9���9�[�9�#�9�(�9�]�9o��9z��9s��9���9[�9`��9�@�9�v�9�=�9[��9�[�9���9���9��9#��9�_�9l(�9"�9Y\�9c��9��9��9x   x   ��9��9�^�9��9�%�9���9*��9�9�+�9�1�9��9k��9v��9;��9�Q�9kS�9b��96��9���9��9�3�9�-�9/�9(��9���9�&�9	��9J_�9���9�9x   x   +��9�^�9�M�9e��9�.�9���9���9���9|��9Y��9H;�9A��9`��9�<�9�t�9;;�9��9��9�;�9{��9���9R��9z��9���9#-�9~��9 N�9C_�9���9ɘ�9x   x   ���9��9F��9���92|�9�*�9���9���9�}�9w�9r�9��9�E�9���9���9�F�9���9kp�9h�9�9��9���9@+�9}�9G��9Ȟ�9C��9 ��9ֈ�9k��9x   x   p[�9a%�9x.�9|�9��9�|�9��9��9�*�9���9˕�9Ur�9���9�"�98��9�p�9|��9S��9�(�9��9��9�{�9���9/|�9�,�9�&�9Q\�9���9���9��9x   x   V#�9t��9���9�*�9�|�9��9oJ�96��9��9~��9��9[n�9s��9N��9Oo�9"��9���9���9N��9�H�9���9*~�9�)�9���9%��94"�9H��9M�9�K�9ߚ�9x   x   X(�9���9f��9z��9��9WJ�9y�93��9M��9�e�9�	�9$a�9k��9�a�9z�91f�9���9���9�y�9�I�9%�9���9F��9���9�(�9�9�:�9 �9�;�9Η�9x   x   �\�9�9}��9���9���9��9'��9%j�9�!�9���9��9d[�9}[�9��9��9w"�9�i�9���9��9[��9i��9���9�9�\�9J��9�t�9M�9�M�9�t�9���9x   x   ���9!+�9���9;}�9�*�9���91��9�!�9}��9��9�@�9�[�9,@�9��9��9 !�9g��9i��9z(�9}�9*��9�,�9&��9�.�9���9i��9��9=��9���9�/�9x   x   ���951�9Ԝ�9�9M��9M��9�e�9��9��9@C�9_U�9V�9_B�9!�9���94d�95��9˄�9��99��9$2�9���9���9�M�9�)�9��9��9�*�9�K�9���9x   x   ���9��9�:�9�q�9|��9���9�	�9��9�@�9`U�9LQ�9�U�9�A�9��9��9v��9V��9mp�9_9�9*�9���9���9���9X��9֧�9H��9���9���91��9���9x   x   ���9ɱ�9���9x��9r�9*n�9a�9S[�9�[�9V�9�U�9�Z�9{[�9�a�9�n�9�q�9���9��9=��9��9���9]�9|�9�)�9�.�9�/�9**�9��9�
�9���9x   x   fZ�9���9��9BE�9���9N��9X��9[�9B@�9iB�9�A�9�[�9P��9���9W��9�F�9���9_��9\�9��9|�9GS�9��9;��9���9���9��9�R�9��9���9x   x   ���9���9<�9;��9�"�94��9�a�9��9��9?�9��9�a�9���9�$�9߫�9k<�9���9ʃ�9&�9v��9�>�9��9���9�9<�9���9���9{=�9���9��9x   x   �?�9ZQ�9Bt�9|��9��9Lo�9��9��9H��9-��9��9�n�9|��9���9�s�9 R�9u?�9"�9���9F��9cg�99��9�:�9 M�9/;�9u��9!h�9���9���9�!�9x   x   [v�9S�9 ;�9bF�9�p�98��9bf�9�"�9E!�9�d�9���9r�9�F�9�<�9R�95u�9���9���9���9���9�v�9�9�B�9�A�9��9�v�9���9���9���9��9x   x   ~=�9"��9ܚ�9���9���9���9��96j�9ʕ�9���9���9\��9ܘ�9E��9�?�9Ģ�9P�9Sa�9��9���9�O�9h��9!��9��9�O�9C��92��9D`�9��9t��9x   x   ��9
��9��9up�9��9���9��9d��9���9H��9�p�9���9���9.��9X"�9��9ma�9���9&!�9��9���9l<�9�;�9���9��9 �9���9�`�9���9 #�9x   x   �[�9��9�;�9��9D)�9���9^z�9l��9)�9�9�9�9��9�\�9��9P��9��9���9C!�99l�9]h�9��9�6�9x�9@i�9�l�9  �9e��9R��9��9��9x   x   ���9��9���9R�9f��92I�9J�9��9�}�9��9��9���9���9��9���9r��9��9  �9}h�9�E�9(��9��9�D�9g�9�!�9���9���9���9,��9j��9x   x   ���9�3�9���9���9�96��9��9%��9���9�2�9i��9���9A�9Z?�9h�9�w�9%P�9���9��9B��9���9s��96�9���9�N�9`y�9�h�9�=�9X�9���9x   x   3��9�-�9���9U��90|�9�~�9���9���9q-�9���9r��9@�9T�9��9���9$�9���9�<�987�9%��9���9B5�9�<�9���9o�9���9��9�T�9�
�9J��9x   x   W��9��9���9�+�9{��9P*�9��9��9	��9��9���9o�9؉�9���9�;�9oC�9���9g<�9��9&E�9a�9�<�9���9C�9�=�9l��9���9z�9*��9$��9x   x   �_�9~��9o��9�}�9�|�9���9���9�]�9y/�9�N�9Y��9�*�93��9�9�M�9�B�9���9C��9�i�9jg�9���9���9C�9�L�9��9���9"+�9,��9�L�970�9x   x   �(�9&��9�-�9���9�-�9���9�)�9:��9���9�*�9ި�90�9���9.�9<�9��9_P�9 �90m�91"�9O�9��9�=�9��9���9'0�9N��9�+�9G��9_��9x   x   X"�9�&�9���9Y��9_'�9�"�9���9�u�9`��9��9V��9�0�9���9���9Y��9�w�9��9!�9z �90��9�y�9��9���9���9)0�9���9�9Z��9u�9��9x   x   �\�9c��9zN�9ڙ�9�\�9��9�;�9�M�9���9��9���9.+�9��9���9�h�9���9ݗ�9=��9ݗ�9���9:i�9>��9��9'+�9Q��9�9:��9^N�9�;�9��9x   x   ���9�_�9�_�9���9W��9�M�9��9�N�9-��9�+�9���9��9�S�9X>�9O��9?��9�`�9a�9���9��9 >�9�T�9~�9*��9�+�9S��9^N�9 �9�L�9,��9x   x   &��9��9[��9I��9���9[L�9L<�9ru�9���9�L�9!��9��9��9f��9V��9T��9�9l��9`��9h��9q�9�
�9&��9�L�9+��9fu�9�;�9�L�9��9���9x   x   �9K�9��9Ј�9���9t��9x��9D��9�0�9W��9���9v��9V��9S �9q"�9���9��9\#�9��9���9���9>��9��90�9,��9��9���9��9���9���9x   x   �o�9С�9$1�9�9�L�9���9�r�9;�9��9���9��9�"�9�d�9]V�9���9�!�9���9�V�9>e�9�"�9ן�9���9��9�<�9�r�9���9TL�9��9q.�9���9x   x   ǡ�9���9;��9a��9Z��9r�9��9��9���95�9���9�
�9��9���9-2�9�3�9w��9�9�
�9B��9�6�9���9���9�9(r�9���9���9]��9* �9��9x   x   �0�9+��9�s�9���9R��9$F�9���9?v�9�	�9���9���9���9���9�N�9�v�9�L�9]��9u��9���9���9��9�v�9���9`E�9F��9��9+r�9��9-/�9O�9x   x   ��9:��9j��9��9���9|=�9���9�(�9���9���9��9P��9G��9���9���9y��9	��9� �9���9K��9�)�9���9�<�9j��9C��9���9���9x�9/��9&��9x   x   NL�9��9��9���9��9�P�9R��9���9t)�9XC�9�*�9���9?@�9Yg�9�?�9��9�+�9�D�9'�9Q��9u��9GP�9��9B��9u��9f��9�K�9���9���9��9x   x   A��9-r�9�E�9Q=�9�P�9�p�9[��9B��9���9K��9M�9���9<�94
�9O��9�M�9���9��9'��9h��9;r�9!Q�9�;�9�F�9_q�9$��9TO�9b�9��9�M�9x   x   r�9h�91��9|��9,��9B��9J��9�t�9?>�92��9�p�9���9x��9+��9*o�9���9�=�90t�9Q��9���9ȣ�98��9���9�9�r�9:��9/��92��9ذ�9���9x   x   �:�9���9�u�9�(�9���9#��9�t�9(�9���9�6�9��9ؿ�9���9��9j7�9���9
(�9Ot�9��9M��9&*�9su�9��9}:�9���9v��9�W�9�X�9��9���9x   x   F�9,��9d	�9M��99)�9̺�9#>�9���9)�96x�9&��9һ�9���9�y�9'�9���9?�9%��9\(�9��9u�9��9�9��9�u�9�E�95=�9�E�9=u�9u��9x   x   ��9�4�9��9���9C�9��9��9�6�94x�9��9���9c��9���9.x�9�9�9���9���9�C�9��9���976�9���9��9{�9T�9�F�9�E�9�U�9�z�9��9x   x   l��9��9e��9@�9�*�9�L�9�p�9��9��9���9-��9���9��9Ԑ�9Nn�9�N�9+�9�9���9���9���9��9�o�9d�9�]�9�[�9�]�9sb�9�p�9��9x   x   �!�9[
�9h��9���9���9���9���9п�9ѻ�9e��9���9r��9Ϳ�9���9��9���9y��9���9v
�9	"�9:�9'L�9&_�9xl�9+v�9Pw�9�l�9n`�9fL�9�7�9x   x   d�9 �9s��9���9	@�9�9f��9���9���9��9 ��9ҿ�9i��9B
�9@�9@��9e��98�9�d�9���9���9T2�9ya�9�u�9���9�s�9�a�9�/�9���9���9x   x   �U�9P��9AN�9���9-g�9#
�9*��9���9�y�9Lx�9��9���9O
�9�g�9���9PM�9���9�U�9���9�Y�9��9�"�9O�9�q�9�r�9�O�9Y$�9���9�V�9V��9x   x   f��9�1�9Fv�9���9�?�9P��9:o�9�7�9)'�9�9�9xn�9B��93@�9���9[v�9�2�9���9��9�_�9���9}��9���9�.�9�J�94.�9���9f��9 �9�a�9���9x   x   �!�9_3�9VL�9^��9��9�M�9���9���9��9���9O�9��9s��9oM�9�2�9� �9F�9��9���9���9|3�9���9���9���9֛�9W4�9ƛ�92��9`�9��9x   x   c��9E��9?��9��9�+�9���9>�9T(�9f?�9��9]+�9���9���9���9���9Y�9�:�9M�9uJ�9�9���9h�940�9��9��9��9bJ�9KL�9�>�9;�9x   x   eV�9d�9p��9� �9 E�98��9xt�9�t�9���9_D�9��9
��9��9V�9/��9��9M�9���9���9`�9$��9�8�9�9�9���9�`�9o��9���9�K�9��9o��9x   x   e�9�
�9���9��9S'�9|��9���9���9�(�9���9r��9�
�9He�9G��9%`�9���9�J�9���9a��9re�9���9�
�9���9'f�9���9��9K�9��9�a�9p��9x   x   �"�9J��9Ј�9���9���9ʛ�9.��9���9���9=��9��9�"�9���9Z�9k �9ߜ�9V�95`�9�e�9i�9kt�95u�9j�9�d�9fb�9��9)��9���9CX�9^��9x   x   ���97�9��9�)�9٥�9�r�9Q��9�*�9�9�6�9A��9�:�9I��9���9���9�3�9��9i��9���9{t�9���9�t�9���9���9���9N5�9���9Y��9/��9l9�9x   x   ���9/��9�v�9���9�P�9�Q�9ҳ�9v�9���9H��9ͅ�9�L�93�9�#�9���9��9��99�9�
�9\u�9�t�9#
�9�9�9��9���9N��9�#�9�1�9�K�9���9x   x   �9���9-��9G=�9�9m<�9O��9���9��9��9�p�9�_�99b�9�O�9q/�9F��9�0�9 :�9���9��9���9�9�9�/�9���9/�9�P�9Ab�9a�9r�9+��9x   x   �<�9_�9�E�9���9���95G�9��9A;�9ֹ�9�{�9�d�9Km�9\v�9`r�94K�9{��9}�9��9|f�9�d�9���9��9��9K�9&s�9"u�9mm�9Ec�9�z�9���9x   x   s�9zr�9���9���9	��9r�9�s�9E��9�v�9�T�9�^�9w�9o��9�s�9�.�9t��9y��9,a�9ݘ�9�b�9ɵ�9ٚ�9*/�90s�9��9=x�9�^�9�V�9w�9}��9x   x   ���9N��9~��9��9���9���9���9A��9\F�9�G�9�\�9(x�9�t�9�P�9���9�4�9�9��9k��9�9�5�9i��9�P�9)u�9<x�9T[�9�G�9�D�9r��9u��9x   x   �L�9ά�9�r�9n��9L�9�O�9ޱ�9�X�9>�9�F�9R^�9�m�9Qb�9 %�9��9g��9�J�9��9sK�9n��9(��9$�9Kb�9nm�9�^�9�G�9�>�9lY�9ȯ�9<O�9x   x   ��9���91��9��9��9��9ڛ�9vY�9YF�9vV�9:c�99a�90�9���9� �9���9�L�9[L�9f��9# �9���9�1�9a�9?c�9�V�9zD�9jY�9���9��9���9x   x   �.�9k �9z/�9���9���94�9{��9e��9�u�9�{�9Tq�9$M�9���9�W�9^b�9��9,?�9.�9b�9nX�9F��9�K�9r�9�z�9�v�9P��9���9��9-��9���9x   x   ���94��9��9}��9q��98N�9��9|��9!��9���9˅�9�8�9c��9���9 ��9�9��9���9���9}��9q9�9���9��9f��9X��9L��9O�9���9���9H�9x   x   w�9p��93�9���9���9e�9�d�9���9�h�9@��9�F�9���9S��9�S�99��9E��9���9�S�9���9���9NG�9U��9i�9k��9xe�9�9���9���9'�94��9x   x   Z��9���9,|�9zL�9�V�9���9��9U�9߼�9��9�X�9Ps�9VQ�9���9d0�9<1�9o��9�P�9�s�9�X�9!�9#��9MS�9[��9�9�U�9�M�9}�9.��9���9x   x   �9|�9�,�9��9)�9U@�9���9���9�*�9�f�9�z�9_�9,�9�{�9A��9�y�9��9�_�97{�99f�9�)�9y��9���9#@�9��9`�9�*�9${�9��9���9x   x   ���9TL�9��9I��9F��9A�9bF�9x�9N��9��9���9L�9g��9��9�9,��9�L�9;��9\��9���9Hw�9�F�9a�9���9|��9x�9O�9��9[��9��9x   x   ���9�V�9�9:��9��9a��9X�9m�9�9G��9ط�9�I�9�9���90��9XH�97��9\��9�9��9)�9���9���9���9^�9�S�9���9`��9^h�9���9x   x   �9���9'@�9�9K��9b��9��9���9Ȍ�9�A�9��9�7�9�p�95p�999�9���9�@�9���9���9#��9��9��9��9�?�9%��9��9ث�9bu�9sw�9���9x   x   `d�9���9d��9<F�9B�9���9���9�V�9E��9"��9C��9:.�9g@�9P.�9���9Ӈ�9���9JV�9���9J��9r�9�F�9H��9���9e�9��96��9"��9���9��9x   x   d��9�T�9���9�w�9C�9���9yV�9���9�f�9e��9�9�$�9%�9W�9k��9vg�9?��94W�9���9��9x�95��9�U�9���9*~�9�F�9~ �9!�9F�9r~�9x   x   h�9y��9O*�9��9��9���9;��9�f�9���9���9��9� �9��9���9Q��9Ef�9���9΍�9
�9��9K+�9Ի�9g�9l�9���9@��9S��9���9���9��9x   x   ���9/�9Xf�9���9��9�A�9��9[��9���9�9�$�9�%�9#�9z��9+��9��9I@�9I��9k��9�d�9s�9��9}��9��9fh�9�b�9�_�9�i�9ކ�9U��9x   x   F�9�X�9�z�93��9���9���9+��9��9��9�$�96.�9�$�9t�9�9o��9���9:��9T��9w{�9�W�9�D�9�1�9�&�9��9��9��9�9F�9B&�9�1�9x   x   !��9�r�9�^�9�K�9\I�9�7�9.�9�$�9� �9�%�9�$�9� �9�$�9�0�9�7�9�F�9DL�9�]�9t�9>��9ӝ�9��9R��9���9���9n��9���9��91��9���9x   x   ڍ�9�P�9��9-��9���9�p�9Y@�9%�9��92�9{�9�$�9u>�90p�90��9���9��9�O�9��9���9��9�4�9~V�9�o�9�t�9n�9aW�9]1�9��9���9x   x   dS�9|��9a{�9��9���9'p�9H.�9c�9���9���90�9�0�9<p�9o��9��9$y�9���90U�9)��91"�9�z�9O��9��9�	�9)�9���9;��9�|�92!�9=��9x   x   ���90�9��9��9��959�9��9���9h��9O��9���9�7�9E��9��9���9p0�9���9i�9 ��9ŀ�9���9\:�9�t�9[��93t�9p8�9&��9=�9���9*j�9x   x   ���9�0�9�y�9��9PH�9���9��9�g�9pf�9E��9���9�F�9���9Ey�9�0�9���9J��9��9[4�9���94G�9��9���9���9���9�H�9���9�5�9=��9M��9x   x   ���9A��9��9�L�9G��9A�9���9y��9���9�@�9���9~L�9+�9���9��9f��9��9#��9NU�9b��9)��9-��9`��9:��9�~�9��9�T�9���9۬�9��9x   x   VS�9iP�9�_�9D��9y��9���9�V�9�W�9��9���9���9I^�9�O�9qU�9Hi�9���9:��9ً�9�]�98�9y��9u��9c��9���9��9^�9 ��9X��9���9�j�9x   x   y��9�s�9C{�9r��9K�9���9֓�9W��9j�9а�9�{�9kt�9ތ�9���9d��9�4�9|U�9�]�9�9�9���9�D�9>c�9QB�9���9�7�9�]�9�U�9�5�9{��9.��9x   x   ���9�X�9Sf�9���9�9y��9���9��9|��9ee�9)X�9���9$��9�"�9#��9���9���9Y�9���9o�9���9���9vp�9b��9��9&��9���9_��9� �9	��9x   x   XG�9;�9 *�9�w�9z�9���9��9�x�9�+�9��9ZE�9]��9�9!{�9/��9�G�9v��9���9 E�9���9���9���9<C�9���9��9?H�9���96}�9:�9���9x   x   j��9O��9���9DG�9X��9{��9"G�9���9i��9���902�9|��95�9ջ�9�:�9���9���9���9uc�9��9���9Wd�9���9���9қ�9�:�9��9�2�9Ȫ�9R3�9x   x   (i�9}S�9��9��9���9�9Ή�9�V�9�g�9��9�'�9��9W�9���9�u�9:��9���9���9�B�9�p�9WC�9��9���9?��9�s�9���9�X�9e��9'�9���9x   x   ���9���9t@�9���9���9@�9,��9}��9�9���9A�9���9yp�9)
�9��9V��9���9���9��9���9���9���9M��9k��9k�9Nn�9���9��9��9��9x   x   �e�9���9��9���9��9���9�e�9�~�9h��9i�9��92��9�u�9��9�t�9;��9�9+�9 8�9+�9:��9��9�s�9o�9Hu�9���9�9�j�9���9�|�9x   x   5�9�U�9��9��9gT�9+�9G�90G�9���9Mc�9��9��9�n�9>��9
9�9I�9���9o^�9�]�9g��9kH�9�:�9���9Wn�9���9��9nb�9���9�I�9Z�9x   x   ���9�M�9�*�9jO�9,��9]��9���9 !�9��9T`�9��9i��9X�9Լ�9���9^��9U�9{��9�U�9���9���9.��9�X�9��9�9ub�9��9g!�9/��9���9x   x   ��9L}�9o{�9o��9ʃ�9�u�9���9�!�9i��9rj�9��9���9�1�9�}�9��96�9`��9���9�5�9���9Q}�9�2�9n��9��9�j�9���9Z!�9��9�w�9��9x   x   C�9O��9��9���9�h�9�w�9��9�F�9"��9}��9�&�9ͫ�9B�9�!�9��9���99��9ʀ�9���9� �9S�9Ϫ�9'�9߅�9���9�I�9��9�w�9�f�9s��9x   x   B��9���9���9^��9���9��9��9�~�9S�9��9c2�9H��9J��9���9�j�9���9b��9�j�9W��9��9���9D3�9���9��9�|�9<�9ի�9���9d��9��9x   x   ��9K:�9G��9q7�9�9��9!�9v]�9���9���9.��9���9���9�o�9���9���9*��9No�9_��9���9\��9���9���9�]�9<"�9��9s�9�6�9���9):�9x   x   <:�9�s�9���9>��9}z�9�u�9��9۹�9���9�9��9���9���9��9�R�9_R�9��93��9��9�9��9���9\��9ˍ�9#s�95z�9M��9���9�t�9�8�9x   x   *��9���9�x�9G(�9��9/�9�9�(�9�8�9�3�9��9���9�a�9g��9���9J��9�a�9s��9��9�2�9�9�9�)�9i�9��9�	�9}(�9fv�9���9ӛ�9Y|�9x   x   N7�9!��98(�9k��9���9��9���9Ĥ�9-��9q�99�9w��9�1�9�k�9dl�9�1�9��9�8�9�q�9��9Ģ�9���9���9S��9X��9�(�9���9�5�9��9w�9x   x   �
�9Lz�9c�9���9���9_�9�B�9O$�9���9g��9_E�9ζ�9��9Y�9s�9���9E�9���9���9�$�9�C�9>`�9z��9\��9�
�9w�9�	�9���9��9��9x   x   N�9zu�9�9ī�9�^�9P*�9���97��99V�9���9`\�9%��9���9���9е�9@\�9���9�V�9U��9���9�'�9�^�9��9�9�u�9�9���9��9���9W��9x   x   � �9̌�9��9���9iB�9���9-��9�(�9˲�9�$�9fy�9��9���9���9�x�9�%�9ͱ�9�(�9���94��9�C�9S��9��9G��9�!�9K��9ˢ�9֓�9v��9<��9x   x   ]�9���9c(�9���9,$�9$��9�(�9	��91��9ZR�9݂�9g��9���9���9�Q�9o��9���9�(�9@��97#�9��94'�9h��9�\�9�9���9)��94��9���9 �9x   x   O��9h��9�8�9���9���9V�9���9&��9�E�9�y�9v��9F��9k��9Dz�9jE�9���9��9�W�96��9��9�:�9���9ƕ�9�Y�9�.�9��9X�9��9�,�9Y�9x   x   n��9��9�3�9�p�9;��9���9�$�9NR�9�y�9q��9ڡ�9��9��9�y�9rR�9�%�9���9ӭ�9�q�9{1�9��90��9���9�~�9�j�9uZ�9W�9k�9���9��9x   x   ���9-�9��9�8�92E�9B\�9Ry�9ق�9w��9ۡ�90��9��9Ɩ�9���9�x�9�\�9xF�9�8�9��9~�9w��9���9���90��9���9��9��9���9���9���9x   x   J��9V��9e��9<��9���9��9���9]��9?��9��9ס�9`��9<��9��9}��9H��9���9~��9���9���9o�9��9~�9'�9(+�9+�9�%�9`�9��9u�9x   x   b��9���9�a�9�1�9��9���9}��9ë�9u��9���9Җ�9E��9ھ�9���9��9�0�9�c�9���9���9X��90�9�T�9�l�9���9���9R��9�m�9GR�9�/�9���9x   x   �o�9��9)��9�k�97�9���9���9���9Tz�9�y�9���9��9���9��9�k�9���9�9q�9d��9>�9�`�9]��9*��9���9���90��9f��9"c�9��9���9x   x   ���9�R�9���9Bl�9c�9е�9�x�9�Q�9�E�9�R�9�x�9���9��9�k�9���9�Q�9���9�O�9!��9�0�9V��9w��9���9���9��9���9��9.�9/��9�P�9x   x   ���94R�9*��9�1�9���9R\�9�%�9���9!��9�%�9]�9t��91�9���9R�9r��9���9�3�9���9�C�9���9��9��9��9���9��9dE�9 ��9�1�9A��9x   x   ���9d�9�a�9���9#E�9���9��9���9��9��9�F�9���9�c�91�9���9��9�T�9T�9ĳ�9�=�9��9V��93��99��9%��9�<�9e��9k�9�U�9E��9x   x   *o�9"��9p��9�8�9���9W�9�(�9�(�9�W�9��9�8�9���9��9Hq�9P�9�3�9b�9���9��9�9r�9���9Q��9�r�9��9��9'��9��92�9�P�9x   x   J��9
��9��9�q�9���9���9��9���9���9r�9 �9M��9��9���9_��9���9޳�9���91>�9���9��9�&�9e�9���9a<�9M��9���9���9p��9���9x   x   ���9�9
3�9.��9�$�9���9���9�#�9u��9�1�9��9���9���9��9>1�9�C�9&>�90�9���9�3�9ws�9ks�9�5�9>��9I�9�>�9D�90�9�9���9x   x   b��9��9�9�9��9D�95(�9'D�9K��9V;�9��9���9��9�0�9a�9���9��9M��9=r�9�9�s�9n��9As�9��9�r�9��9��9r��9�c�9]1�9� �9x   x   ���9���9�)�9ߢ�9�`�9B_�9���9�'�9��9���9(��9�9"U�9ǔ�9���9p��9���9��9�&�9�s�9Is�9�(�9��9���9?��9m��9���9�R�9��9���9x   x   ݗ�9���9��9۪�9҉�9Q��91�9��9F��9��9y��9��9<m�9���99��97�9���9���9��9#6�9��9��9���9��9���9%��9�n�9=�9I��9X��9x   x   �]�9���9��9���9���9��9���9[]�9NZ�9"�9���9�'�9E��9]��9`��9/�9���9�r�9ھ�9n��9�r�9���9��9I��9���9߅�9�&�9���9��9cY�9x   x   i"�9Vs�92
�9���9!�92v�9R"�9��9F/�9}k�9S��9�+�94��95��9���9���9��9��9�<�9w�9C��9T��9���9���9���9�,�9=��9�l�9�.�9��9x   x   &�9fz�9�(�9)�9nw�9y�9���9N��97�9 [�9���9�+�9݆�9���9u��9_��9.=�9A��9���9?�9��9���92��9ޅ�9�,�9���9�Y�9h�9���9���9x   x   ��9���9�v�9��9X
�9��9C��9���9��9�W�9���9w&�9'n�9��9^��9�E�9���9x��9���9,D�9���9���9�n�9�&�97��9�Y�9s�9,��9?��9o��9x   x   �6�9���9��96�9���9��9K��9���9x�9�k�9��9��9�R�9�c�9z.�9g��9��9��9$��990�9�c�9�R�9@�9���9�l�9]�9)��9T��9h��9h��9x   x   ��9 u�9��9�9k��9
��9��9q��9j-�9>��9��9�9T0�9Y�9���9I2�9V�9U2�9���9$�9r1�9��9D��9��9�.�9���92��9[��9��9��9x   x   6:�9�8�9|�9��9d��9���9���9k�9�Y�9���9c��9��9d��9���9Q�9���9���9�P�9���9���9� �9���9K��9JY�9��9���9U��9R��9��9�|�9x   x   @b�9�u�9���9�C�9{��9���9��9ʡ�9J��9��9��9Yo�9"�9���9���9Z�9O��9V��9�9'n�9��9��9Φ�9��9;��9ֻ�9@��9cB�9���9�u�9x   x   �u�9Z��98�9.��9�L�9��9<�9?��9���9r��9ǩ�9�_�9���9�\�9���9���9R\�9a��9
`�9S��9���9Z��9���9��9$�9M�9���9��9���9�r�9x   x   ���9(�9�y�9��9J��94��9q�9zP�9�,�9~ �9	��9Q�9���9�
�9� �9J�95��9�O�9��9���9�-�9�Q�9�r�9ܔ�9-��9+�9Vw�9��9���9ܯ�9x   x   wC�9��9��97��9�T�9��9B��9��9v{�9�0�9��9I�9���9U��9,��9���9�I�9���9�0�9�{�9��9R��92�9�U�9���9;�9
��9-@�9�9��9x   x   G��9pL�90��9�T�9���9���9Wn�9�&�9\��9f�9W��9g=�9�w�9���9�w�9L>�9���9Ve�95��9G'�9(p�9���9���9T�9���9!J�9���9#��9W��9ж�9x   x   e��9��9��9��9���9|O�9O��9���98�9���9���9�5�9�V�9�W�9�5�9���9���9�9{��9v��9�M�9ͺ�9�9��9H�94��9m��9-c�9ld�9�9x   x   ή�9
�9�p�9&��9An�9C��9�u�9��9�e�9���9��92-�9�<�9I,�9i�9
��9�c�9���9�v�9"��9lo�9H��9tq�9��9i��9�n�9?�9�/�9R?�9Oo�9x   x   z��9
��9GP�9ζ�9k&�9���9��9X�9���9}��9?�9�(�9&)�9�9��9���9�X�9���9���9�%�9���9kP�9���9��9�m�9�9�9`(�9�'�9�8�9In�9x   x   ���9���9�,�9K{�93��9$�9�e�9~��9��9��9��9"�94�9��9���9٩�9~e�97�9���98{�9�-�9��9���9�w�9pQ�9�7�9�5�9�9�9TQ�9�v�9x   x   Ī�9(��9< �9�0�9�e�9���9���9z��9��9��9<&�9
'�9��94�9���9��9N��9Qd�91�9O��9���9x��9V��9�l�9S[�9�U�9hS�9ZZ�9_m�9���9x   x   ���9{��9ɷ�9���93��9��9��9;�9��9=&�9i,�90&�9t�9��9	�9���9X��9���9���9F��9���9���9Ά�9�{�9�x�9xx�9�{�9-{�91��9��9x   x   �n�99_�9�P�9�H�9J=�9�5�9!-�9�(�9"�9'�92&�9�"�9(�9�+�9�4�9�=�99I�9(O�9�`�9�m�9�{�90��9P��9�9;��9���9Ҕ�9w��9>��9�{�9x   x   ��9l��9z��9^��9�w�9�V�9�<�9)�96�9��9~�9�(�9E>�9�V�9y�9���9���9���9��9�J�9Sd�9;��9N��9���9Ϻ�9���9J��9ٌ�9Ld�9�I�9x   x   <��9�\�9�
�97��9���9}W�9K,�9�9��9?�9��9�+�9�V�9���9&��9j�9$\�9L��9���9�.�9�`�9��9��9���9���9���9֛�9,b�9�/�9���9x   x   g��9L��9` �9��9�w�9�5�9q�9)��9���9���9$�9�4�9y�9.��9!�9���9���9�X�9��9$�9�]�9ŏ�9��9���9���9���9�]�9��96��9�X�9x   x   �9���9(�9���9G>�9���9��9ͩ�9���9���9���9>�9Ş�9y�9���9�9��9�9|��9'��9�=�9�v�9���9��9Ev�9<�9��9���9��9G��9x   x   '��93\�9#��9�I�9���9���9d�9�X�9�e�9q��9���9eI�9���9I\�9��9��9�5�9���9�M�9 ��9�	�9�B�9O�9�A�9��9��9�K�9���9�5�9���9x   x   =��9S��9�O�9���9he�97�9���9���9j�9�d�9���9aO�9���9~��9�X�9!�9���9�g�9Z��9�i�9R��9��9���9��9�j�97��9�h�9��9�9�X�9x   x   ��9 `�9��9�0�9S��9���9w�9��9$��9R1�98��9�`�9��9���9��9���9�M�9e��9�~�9$��97�9�R�9�7�9���9�~�9���9K�9و�9���9��9x   x   !n�9U��9���9
|�9r'�9���9b��9&�9�{�9���9���9�m�9BK�9�.�9Y�9X��9F��9j�94��9�N�9%��9���9�P�9���9^h�9x��9#��9��9[-�92L�9x   x   "��9���9.�98��9_p�9�M�9�o�9ж�9.�9��9��9|�9�d�9�`�9 ^�9�=�9)
�9v��947�94��9S��9��94�9���9�	�9�<�9�]�9)c�9�d�9�{�9x   x   ��9y��9�Q�9���9��9��9���9�P�9k��9��9��9���9���9u��9��9�v�9C�9F��9S�9���9��9bU�9���9C�9�v�9���9���9'��9��9Г�9x   x   ��9���9�r�9j�9C �9T�9�q�9��9��9���9<��9���9���9w��9i��9��9^O�9��9�7�9�P�914�9���9�M�9M��9Э�9Ѭ�9���9���9��99��9x   x   ��9�9��9V�9QT�9H��9`�9v��9x�9�l�9|�94��9��9���9S��9:��9�A�9$��9���9 ��9���9C�9R��9L��9y��9���9*��9!{�9�m�9�v�9x   x   W��9S�9c��95��9K��9��9ɰ�9n�9�Q�9�[�9Qy�9���9B��9I��9��9�v�9�9�j�9�~�9�h�9�	�9�v�9߭�9���9{��9v��9�z�9\�9�Q�9dn�9x   x   ��9=M�9j�9��9rJ�9���9o�9$:�928�9BV�9�x�99��9���9���9O��9a<�97��9x��9���9���9�<�9���9Ҭ�9���9���9jx�9�T�9�7�9$;�9m�9x   x   ]��9٘�9�w�9I��9B��9Ā�9�?�9�(�9C6�9�S�9|�9H��9���9?��9�]�9v��9;L�9i�9PK�9Q��9�]�9���9���9(��9�z�9�T�9I8�9�'�9o@�9���9x   x   yB�9��9��9e@�9o��9c�90�9P(�9 :�9�Z�9�{�9��9F��9�b�91�9��9���98��9���9�9?c�98��9Ē�9!{�9\�9�7�9�'�9l0�9�c�96��9x   x   ���9���9���9E�9���9�d�9�?�9�8�9�Q�9�m�9���9���9�d�9�/�9���9��9�5�9;�9���9s-�9�d�9���9؆�9�m�9�Q�9;�9d@�9�c�9#��9c�9x   x   �u�9�r�9���9)�9��9��9�o�9�n�90w�9��9D��9M|�9AJ�9=��9 Y�9���9��9�X�9=��9?L�9�{�9Γ�9*��9�v�9On�9�l�9{��9*��9]�9���9x   x   �Z�9�k�9���9~�9ߨ�9�K�9;�9O��9c��9�}�9�?�9���9��9 ��9b+�9?@�9I-�93��9�~�9I��9�@�9h~�9���9T��9+�9M�9	��9�9���9l�9x   x   �k�9`��91��9zX�9I��9͗�9'V�9��9��9i��9dL�96��9W_�9���9A��9d��96��9�a�9���91L�9��9d��9��9V�9R��9P��9�Z�9���9���9_j�9x   x   o��9'��9\B�9!��9�J�9���90��9�d�9��9T��9�b�9���9�7�9os�9b��94u�9W7�9���9c�9���9��9�e�9��9R��9yJ�9.��9QA�9���9`��9��9x   x   a�9cX�9��9�9�9���9�f�9��9��9�Z�9q��9|e�9���9�9[<�9�;�9�9���9g�9���9TZ�9ǵ�9��9ze�9���9�:�9B��9mY�9;�9���9���9x   x   ���9+��9�J�9���9HO�9R��9�z�9Y
�9O��9��9U|�9���9	��9I�9���9���9Y{�9��9m��9Y�9({�9���9[P�9���9oJ�9���9��9�w�9�^�9�u�9x   x   zK�9���9���9zf�9F��9#e�9w��97i�9���9 :�9���9¿�9���9���9N��9J��9m;�9f��9*g�9'��9�d�9���9�f�9��9���9<K�9)�9R��9O��9��9x   x   ��9�U�9
��9��9�z�9p��9qZ�9,��9[�9[�9���9ո�9���9 ��9���9\�9��9��9\�9 ��9�{�9��9��98V�9{�9���9\��9���9&��9��9x   x   ��9��9�d�9ƶ�9?
�9+i�9#��9��9	I�9�~�9b��9��9-��9���9v}�9�H�9��9��9�h�9�	�9׶�9�e�9��9%��9���9���9Oy�9�x�9/��9���9x   x    ��9���9��9�Z�98��9���9L�9�H�9 m�9ݗ�9���9���9X��9���9(n�9�I�9��9���9���9\Z�9x�9���9ڷ�9l��9�i�9�W�9�M�9�X�9/j�9*��9x   x   ^}�94��9$��9K��9��9�9�9[�9�~�9֗�9-��93��9��9��9L��9�|�9VZ�97<�9��9���9���9���9�|�9�`�9�L�9�>�9{7�9R6�9f=�9 M�9b�9x   x   �?�9-L�9�b�9Ue�97|�9���9���9^��9��9(��9��9��9���9<��9���9k��9�{�9g�9�a�9@L�9�@�9�2�9.)�9�)�9��9��9%"�9s*�9'�9d3�9x   x   ���9��9���9���9s��9���9˸�9��9���9���9��9���9���99��9:��9��9���9���9w��9Z��9$��9Z�9
�9%�9<�9�9��9��9f�9J��9x   x   ��9&_�9�7�9��9���9���9���9*��9U��9��9��9���9}��9��9g��98�9~7�9�`�9��9s��9���9���9?��9e��9��9���9���9���9I��9 ��9x   x   ���9Ĭ�9Js�9<<�99�9���9���9���9�9X��9I��9@��9��9��9<�9pu�9ޫ�9���9"�9p[�9���9@��9���9��9#��9���9��9ʈ�9P\�9� �9x   x   ,+�9 ��9?��9�;�9���9G��9���9�}�9<n�9�|�9̙�9G��9u��9<�9���9���9�-�9���9���9�9iS�9ހ�9w��9��9ߛ�9��9S�9��9���9���9x   x   @�9I��9%u�9��9���9P��9\�9�H�9�I�9nZ�9���9+��9P�9�u�9���96@�9���9;�9Sy�9,��91�9�@�9�N�9WP�9�>�9��9���9y�9��9S��9x   x   $-�9��9K7�9���9g{�9~;�9��9��9��9c<�9�{�9	��9�7�9���9�-�9���9�+�9S��9��9}o�9õ�9��9���9���9͸�9�n�9Z�9��9�*�9K��9x   x   ��9�a�9���9g�9��9~��9&��9��9���9��9Jg�9���9�`�9���9���9J�9\��9�5�9���9
�9n;�9�\�9�\�9�:�9-�9���9�6�9��9J�9���9x   x   �~�9���9"c�9���9���9Rg�92\�9i�9ݚ�9*��97b�9���9-��99"�9���9py�9��9���9��9�q�9���9��9���9Dp�9D�9֨�9��9	z�9_��9�"�9x   x   E��98L�9���9hZ�9{�9T��98��9�	�9�Z�9+��9�L�9���9���9�[�9M�9R��9�o�9�9�q�9���9���94��9<��9�r�93 �9�q�9���9n�9�Z�9���9x   x   �@�9���9	�9��9T{�9e�9|�9��9��9��9&A�9l��9���9���9�S�9\�9��9�;�9���9��9���9���9���9�<�9۶�9��9�R�9ۉ�9i��9M��9x   x   p~�9w��9�e�9��9���9���9�9f�9���98}�9L3�9��9���9���9!��9�@�94��9�\�96��9B��9���9���9]�9���9�?�9���9��9���9�9�2�9x   x   ���9��9-��9�e�9�P�9$g�9g��9�9.��9.a�9�)�9y
�9���91��9ě�9�N�9��9]�9���9W��9���9
]�9��9oP�9���9���9��98�9�)�9�`�9x   x   q��9(V�9}��9���9���9Y��9�V�9~��9̈�9>M�9G*�9��9���9Y��9:��9�P�9��9;�9lp�9�r�9�<�9���9oP�9M��9��9K��9��93)�9ON�9��9x   x   D�9q��9�J�9;�9�J�9��9��9 ��9j�90?�9 �9��9��9x��90��9G?�9��9^�9q�9U �9��9�?�9���9��9��9_�9""�9�>�9�i�9���9x   x   2M�9o��9Y��9x��9���9�K�9W��9݋�9�W�9�7�9 �9k�9���9��9`��97�9o�9���9���9r�9��9���9���9I��9^�9��9�6�9�X�9B��9���9x   x   #��9�Z�9�A�9�Y�9Q��9k�9���9�y�9N�9�6�9�"�9L�9>��9J��9fS�92��9��97�9��9���9�R�9��9��9��9"�9�6�94O�9�x�9K��9��9x   x   1�9��9���9q�9x�9���9ߨ�91y�9
Y�9�=�9�*�93�94��9��9�9�y�9V��9��9,z�9��9��9���9>�93)�9�>�9�X�9�x�9~��9[��9ax�9x   x   ���9Ɛ�9���9���9_�9���9l��9���9�j�9tM�9�'�9��9���9�\�9��9�9�*�9w�9���9�Z�9w��9�9�)�9@N�9�i�97��9>��9W��9�^�9���9x   x   l�9oj�9@��9���9�u�9��9S��9Ȥ�9r��9Qb�9�3�9���9H��9=!�98��9���9n��9���9�"�9���9T��9�2�9�`�9��9���9���9��9Qx�9���9��9x   x   ��9�&�9�Z�9���9\�9���9CK�9��9���9�M�9��9�|�9���9[L�9�~�9��9��9jJ�9���9"}�9A��9O�9Ҟ�94��9J�9J��9��9���9A]�9�&�9x   x   �&�9	K�9S��9���9�`�9���9���9�$�9���9�j�9���9em�9���9��9�8�9�7�9n�9���9�m�9���9�i�9)��9o%�9��9���9�_�9P��9��9�I�9-(�9x   x   �Z�9M��9���9�6�9��9Z=�9j��9�f�9X��9��9|��9<i�9O��9���9���9���9[��9Hg�9w��9��9���9Wf�9���9d=�9T��9�5�9���9���9�Y�9/I�9x   x   ���9���9�6�9P��9"�9��9o!�9���9�,�9���9��9=b�9K��9-��9c��9s��9�b�9��9<��9�*�9��9�"�9[��9��9���9�5�9��9d��9��9���9x   x   ?�9�`�9m��9�9Z��9���9�w�9���9�_�9���9��9�S�9��9}��9�9�T�9x�9w��9;b�9���9Iv�9��9���9?�9���9b�9��9���9���9}��9x   x   s��9���9E=�9ښ�9���9�k�9���9�6�9ٖ�9��9�"�9DS�9Vf�9�f�9�R�9�!�9���9͖�9�4�9���9�l�9��9ě�9%=�9���9ձ�9�}�9&o�9kp�9�}�9x   x    K�9˃�9T��9[!�9�w�9���9"�9�{�9A��9��99.�9�L�9%Y�9nL�9�.�9��9`��9|�9�"�95��9#y�9� �9���9p��9�I�9�9��9k��9��94�9x   x   ���9z$�9�f�9۫�9���9�6�9�{�9��9���9��9�.�9"G�9G�9	/�9!�9���9ʹ�9�{�9�6�9��9���9<g�97#�9i��9k��9p��9Ý�9���9��9���9x   x   r��9���96��9�,�9�_�9ʖ�9<��9���9r�9�.�9�<�9uH�9�<�97.�9��9���9���9��9�a�9(,�9���9���9���9��9�f�9>T�9�K�9�T�9�f�9��9x   x   �M�9�j�9��9]��9���9n��9x�9��9�.�9>>�9�E�9�E�9l>�9�.�9��9��9p��9���9��9A��9Qi�9N�9$5�9�#�9c�9�9�9�9�$�95�9x   x   D��9x��9R��9��9��9�"�91.�9�.�9�<�9�E�9�E�9�E�9�<�9�/�9�/�9: �9��9��9���9N��9���9w��9��9I��9���9V��9q��9���9���9���9x   x   d|�91m�9i�9!b�9�S�9:S�9�L�9G�9uH�9�E�9�E�9�H�9�F�9K�9�S�9MU�9�a�9�g�9m�9,}�9�~�9���9؏�9���9���9Ƙ�9��9:��9���9h�9x   x   ���9���9*��9-��9��9Jf�9Y�9G�9�<�9s>�9�<�9�F�9�Z�96f�9�~�9���9���9���9���9��9q&�9�<�9�C�9DP�9mK�9�R�98D�9�<�9�$�9q�9x   x   *L�9��9���9��9q��9�f�9kL�9/�9@.�9�.�9�/�9K�9>f�9:��9*��9��9��9�J�9�z�9>��9���9���9)�9(�9��9��9���9���9��97y�9x   x   r~�98�9���9N��9v�9�R�9�.�9*�9��9��9�/�9�S�9�~�9-��9��98�9��9���9]�9�:�9=j�9��9��9(��9���9"��9mi�9C:�9��9���9x   x   ��9�7�9���9e��9�T�9�!�9
�9���9���9��9O �9iU�9���9��98�9ߒ�9N��9K>�94��9���9��9�&�9�;�9�<�9�$�9��9��9J��94?�9j��9x   x   ��9Y�9R��9�b�9y�9���9r��9��9���9���9��9�a�9��9��9��9Z��92S�9���95
�9ET�9C��9���9���9��93��9{T�9G
�9���9�Q�9���9x   x   YJ�9���9Dg�9��9���9���9>|�9�{�9$��9���9�9�g�9���9�J�9���9]>�9ʷ�9�9�{�9m��98��9\�9k�9���9���9�z�9��9��9�?�9���9x   x   ���9�m�9~��9J��9Sb�9�4�9�"�97�9�a�9N��9��9/m�9���9�z�9{�9G��9B
�9�{�9���9$�9�R�9n^�9�R�9>#�9v��9L|�9��9���9��9H{�9x   x   }�9���9���9�*�9���9���9Z��9F��9Z,�9v��9���9Y}�9��9m��9;�9���9_T�9���9 $�9c�9���9��9cd�9�#�9���9JU�9���9;�9b��9#�9x   x   I��9�i�9���9���9rv�9�l�9Oy�9ث�9��9�i�9���93�9�&�9��9nj�9��9f��9S��9�R�9���9:��9~��9�Q�9`��9���9��96i�9T��9�%�9,�9x   x   O�9?��9tf�9�"�9A��9G��9.!�9ug�9���9aN�9���9=��9,=�9���9A��9'�9ŭ�9|�9�^�9��9���9�^�9��9B��9-&�9��9��9�<�9��9���9x   x   ��9�%�9��9���9���9���9 ��9z#�9A��9l5�9R��9��9=D�9k�9=��9�;�9��9��9�R�9wd�9R�9��9W��9�<�9˦�9"�9E�9n��9���9L4�9x   x   M��96��9�=�9�9r�9a=�9���9���9��9C$�9���9���9�P�9q�9e��9�<�9C��9���9\#�9�#�9q��9T��9�<�9���9��9�Q�9��9���9(&�9M��9x   x   J�9��9|��9���9۰�9���9J�9���98g�9��9��9��9�K�9��9.��95%�9m��9��9���9���9���9:&�9˦�9��9L�9���9���9��9�e�9e��9x   x   b��9
`�9�5�9 6�9Ab�9��9E�9���9�T�9��9���9��9ES�9��9e��9��9�T�9{�9p|�9jU�9��9"��9(�9�Q�9���9���9��9�U�9��9��9x   x   ��9i��9���9<��9��9�}�9��9��9�K�9Z�9���9b��9�D�9F��9�i�9A��9y
�9��9��9���9Ei�9��9E�9��9���9��9L�9@��9�9�}�9x   x   ���9��9���9���9���9`o�9���9̝�9	U�9c�9:��9|��9?=�93��9�:�9z��9��9���9Ɍ�9-;�9b��9�<�9q��9���9��9�U�9<��9���9�o�9P��9x   x   M]�9�I�9�Y�9D��9��9�p�9��9_��9g�9%�9��9��9%�9��9.�9f?�9�Q�9�?�9��9o��9�%�9��9���9%&�9�e�9��9�9�o�9Y��9���9x   x   �&�9>(�9AI�9���9���9�}�9l�9���9#��9\5�99��9��9��9ky�9��9���9��9���9R{�9)�9+�9���9F4�9E��9[��9��9�}�9H��9���97G�9x   x   ��9��9���9v"�9�}�9=��9�o�9[��9	��9(�9@��9�	�9Dj�9��9z��9Y��9���9ެ�9j�9,�94��9��9ƈ�9i��9�n�9���9t~�9�!�9���9(��9x   x   ��9���9��9M�9���9��9���9M(�9��9�)�9���9�9�Q�9���9���9���9d��9eR�9/�9���9d(�9ح�9�*�9��9��9���9�M�9���9a��9���9x   x   ���9��9�8�9P��9Q��9Ca�9=��9W�9m��9�C�9���9���9q=�9�a�9�k�9Ua�9<>�9���9A��9�E�9���9�U�9���9a�9���9ݏ�9�9�9l��9E��9_��9x   x   _"�9M�9J��9y��99?�9"��9�9���9���9l_�92��9��9�!�9O:�9M;�9�!�9���9���9^�9���9g��9��9���9�=�9���9t��9~K�9z$�9	�9	�9x   x   �}�9���9G��92?�9���9�92c�9���9l%�9�v�9	��9��9x�9a�9��9���9M��9�u�9�'�9���9�`�9Q�9ϡ�9%?�9���9V��9v{�9_�9�T�9�^�9x   x   ��9��91a�9��9�9�S�9��9�9J�9K��9i��9S��9���9i��9w��9���9��9�I�9��9���9xU�9��9��9�`�9�9���9���9���9"��9���9x   x   �o�9���9!��9�9$c�9��9���9>�9�u�9v��9l��9Q��9���9���9���9'��9�u�9>�9���9:��9�c�9��9���9Ƣ�9n�9VR�9�5�9!-�9�5�9�R�9x   x   .��9*(�9�V�9ދ�9���9��9>�9�p�9J��9���9��9���9���9���9���9}��9�p�9?�9/�9���9d��9dW�9�'�9���9���9K��9h��9���9|��9��9x   x   މ�9���9K��9���9Y%�9J�9�u�9I��9
��9	��9N��9���9���9��9��9ϖ�97t�9�H�9�&�9u��9���96��9\��9�l�9NY�9+N�9P�9�N�9pY�9Hl�9x   x   ��9a)�9�C�9L_�9�v�9B��9i��9���9��9��9K��9���9���9���9���9ޥ�9o��9Yv�9B]�9mE�92(�9��9��9W��9
��9��9��9��9"��9��9x   x   ��9g��9���9��9��9V��9a��9���9K��9S��9���9K��9)��9p��9���9���9���9X��9���9���9��91��9���9/��9��9*|�9=��9`��9���9���9x   x   �	�9��9w��9���9 ��9A��9L��9���9���9���9F��9V��9���9���9���9���9���9{��9��9a�9��9��9z�9H �9< �9I�99 �9��9�9J�9x   x   j�9�Q�9R=�9�!�9l�9���9���9���9���9���9,��9���9���9G��9��9r"�9�=�9	S�93i�9��9ʐ�9��9l��9��9���9��9��9£�9N��9I��9x   x   ­�9y��9�a�99:�9P�9^��9���9���9���9���9x��9���9K��9d�9�:�9Ha�9���9l��9���9=��9e�9�9�9�B�9�T�9�T�9�A�989�9��9���9��9x   x   X��9���9�k�9@;�9��9u��9���9���9��9���9��9���9��9�:�9�j�9b��9���9�9"N�9,w�9���9���9	��9���9>��9���9#��9Fx�9tN�9��9x   x   E��9���9Fa�9�!�9���9���97��9���9��9���9���9���9}"�9Ra�9n��9w��9X3�9�x�9n��9���9�9=�9�N�9O�9�<�9X�9A��9���9�y�9�3�9x   x   ���9R��9.>�9���9M��9��9
v�9�p�9Lt�9���9���9���9�=�9ˍ�9���9\3�9��9���9.'�9`�9���9���9 ��9	��9n��9�`�9N(�9@��9͍�9�1�9x   x   Ӭ�9aR�9���9��9�u�9�I�9!>�9*?�9�H�9�v�9y��9���9&S�9���9�9�x�9���9u6�9��9���9���9���9/��9���9ܼ�9���9�5�9f��9d{�9��9x   x   j�90�9@��9#^�9�'�9��9��9Q�9�&�9h]�9���9��9Qi�9��9:N�9���9<'�9��9���9~�9c0�9�7�9.0�9x�9���9���9�'�9���9fM�9���9x   x   0�9���9�E�9���9���9���9[��9��9���9�E�9Ǟ�9��9��9a��9Kw�9���9,`�9ƽ�9��9�7�9�U�9V�9�7�9��9F��98_�9z��9�w�9���9���9x   x   6��9n(�9���9���9a�9�U�9�c�9���9���9g(�9F��9��9���9��9��9=�9���9 ��9m0�9�U�95m�9�U�9?1�9���9��9h�9���9��9���9&�9x   x   ��9��9�U�9��9q�9��9��9�W�9f��9��9_��9��9��9:�9���9�=�9ˤ�9���9�7�9V�9�U�97�9w��9���9�=�9P��9{9�9��9P�9���9x   x   ֈ�9�*�9���9ƫ�9���9F��9��9�'�9���9�9��9��9���9�B�96��9 O�9@��9J��9C0�9�7�9M1�9t��9���9�N�9c��9nB�9^��9y�9���9��9x   x   u��90��9 a�9>�9L?�9a�9���9���9�l�9���9r��9� �9���9�T�9��9=O�9+��9���9��9��9���9���9�N�9@��9�T�9��9��9���9���9�m�9x   x   �n�9��9���9���9���96�9Un�9���9�Y�9I��9���9| �9-��9�T�9|��9�<�9���9���9���9T��9��9>�9r��9�T�9���9��9���9���9�W�9���9x   x   ���9���9���9���9���9���9�R�9���9jN�9J��9h|�9��9O��9B�9��9��9�`�9ق�9Ȅ�9R_�9x�9T��9qB�9
��9��9`|�9��9�P�9ſ�94S�9x   x   �~�9�M�9�9�9�K�9�{�90��9�5�9���9LP�9J��9v��9t �9!��9k9�9W��9q��9y(�9�5�9(�9���9���99�9d��9��9���9��9�N�98��9�5�9���9x   x   �!�9���9���9�$�9'_�9ߺ�9R-�98��9�N�9F��9���9��9���9'�9zx�9-��9c��9���9۷�9�w�9��9��9y�9���9���9�P�98��9�-�9ֺ�9�^�9x   x   ���9s��9b��92	�9�T�9K��9�5�9���9�Y�9Z��9���9=�9���9��9�N�9�y�9��9y{�9}M�9���9���9T�9���9���9�W�9���9�5�9ͺ�9�U�9 	�9x   x   2��9���9n��9	�9_�9���9�R�9Q��9{l�9!�9���9�9���97��9��9�3�9 2�9��9���9���9'�9���9��9�m�9���9"S�9��9�^�9��9���9x   x   )�9��91�9�k�9޺�92�9��9���9�f�9f��9)B�9���9���9�,�9�P�9Z�9R�9�-�9 ��9a��9�@�9Q��9�d�9"��9��91�9<��9�k�902�9�9x   x   ��9�'�9�R�9W��9���9TB�9k��9�9$��9r��9�I�9���9y��9��9��9��9��9���9���9�H�9���9q��9�9���9B�9���9��9�R�9i&�9�9x   x   1�9�R�9���9z��9.�9=v�9���9=�9���9C��9�Q�9���9���9���9���9 ��92��9��95Q�9���9���9D;�9_��9v�9��9���9���9�S�9�0�9F)�9x   x   �k�9J��9r��9;�9^�9ۮ�9�9�i�9U��9��9HS�96��9$��9���9���9A��9׍�9"T�9!�9߽�9�l�9z�9&��9�]�9��9���9��9�l�9bZ�9�Z�9x   x   ˺�9���9#�9�]�9��9���9�J�9e��9D��9()�9 `�95��9��9u��9x��9w��9n`�9z(�9���9���9�H�9���9��9�^�9��9?��9y��9w��9��9$��9x   x   �9@B�9/v�9Ү�9���99�9ц�9[��9��9DB�9�h�9�|�9j��9��9�|�9gi�9XB�92�97��9p��9�:�9���9:��9�v�9�@�9��9#��9���9���9���9x   x   ��9U��9���9�9�J�9ʆ�9q��9���9'%�9O�9�j�9:|�9n��9�|�9@j�9�M�9R&�9J��9���9���9HI�9�9z��9���9H��9x^�9�N�9WJ�9P�9�^�9x   x   ���9��9=�9�i�9Z��9X��9���9��9�E�9l]�9�x�9;z�9�y�9�w�9Z_�9�E�9"�9���9=��9���9�i�9�=�9�9?��9���9p��9��9`��9]��9l��9x   x   ff�9��9���9?��98��9��9%�9�E�9�V�9�i�9!z�9�z�9�z�9i�9�U�9�E�94%�9��9"��9���9̜�9���9/f�9TO�9S>�9�/�9Z)�90�9�?�9gN�9x   x   ?��9V��9(��9��9)�9;B�9O�9h]�9�i�9�r�9�z�9dy�9ds�9j�9L^�9<O�9�B�9z*�9z�9* �9���9���9m��9���9C��9���9O��9���9g��9���9x   x   B�9�I�9�Q�92S�9`�9�h�9�j�9�x�9z�9�z�9%~�9�z�9ly�9�x�9�i�9mh�9�^�9�T�9�Q�9H�9FB�9";�9�2�9p3�9�5�92�9n5�9+3�9,4�9�:�9x   x   ���9���9���9"��9)��9�|�95|�9>z�9�z�9dy�9�z�9�z�9�z�9|�95~�9���9X��9���9|��9���9���9��9²�9���9���9s��96��9{��9��9ۮ�9x   x   ���9[��9���9��9��9c��9f��9�y�9�z�9hs�9ly�9�z�9 ��9k��9;��9{��9|��9-��9���9s�9��9��9�+�9G,�94�9�*�9�+�9��9��9x�9x   x   �,�9��9���9���9p��9��9�|�9�w�9i�9'j�9�x�9|�9p��9Ӯ�9���9f��9�9�,�9�D�9�f�97~�9��9���9f��9��9v��9���9i}�9!e�9�D�9x   x   �P�9t�9���9���9u��9�|�9Aj�9b_�9�U�9W^�9�i�9;~�9B��9���9���9��9GQ�97��9Ŧ�9f��9t��90�9�9��9��9y�9R��9���9��9z��9x   x   �Y�9��9���9:��9v��9li�9�M�9�E�9�E�9AO�9yh�9��9���9o��9��9CX�9���9���9��9�-�9N�9�n�9�s�9�s�9o�9�N�9U,�9� �9f��9Ø�9x   x   �Q�9��9*��9Ӎ�9q`�9`B�9Y&�96�9J%�9�B�9�^�9l��9���9)�9OQ�9���9���9��9uW�9ۃ�9���9��9���9A��9V��9���9�X�9��9���9;��9x   x   �-�9���9���9(T�9�(�9A�9Y��9���9��9�*�9�T�9���9B��9�,�9L��9���9��9�d�9���9���9���9��9(�9���9���9��9+c�9��9���9�9x   x   ���9���96Q�9-�9���9L��9���9X��9<��9��9�Q�9���9��9�D�9ݦ�9��9�W�9���9���9��9�*�97�9�+�9w�9���9���9`Y�9���92��9'E�9x   x   [��9�H�9���9��9Ȕ�9���9ԅ�9Ė�9���9N �9?H�9���9��9�f�9���9�-�9���9���9��9@�9#P�9�P�9_>�9��9���9��9�.�9���9g�9� �9x   x   �@�9���9���9�l�9�H�9;�9iI�9�i�9���9���9kB�9���9��9a~�9���9N�9���9���9�*�9&P�9cZ�9OP�9�,�9���9��98M�9��9 }�9�9|��9x   x   W��9��9X;�9��9���9���9C�9>�9���9���9R;�9��9��9-��9R�9o�98��9��97�9�P�9NP�9m6�9j�9o��9_p�9��9k��9��9��9u;�9x   x   �d�9#�9k��9=��9��9X��9���9C�9_f�9���9�2�9��9�+�9)��9.�9t�9���9A�9�+�9f>�9�,�9i�9w��9�r�9��96��9�+�9<��9i3�9 ��9x   x   +��9���93v�9�]�9�^�9�v�9"��9i��9�O�9���9�3�9ٴ�9y,�9���9�9�s�9e��9���9��9��9���9y��9�r�9�9���9�,�9���9�4�9;��9�P�9x   x   ���9B�9��9��9��9"A�9w��9���9�>�9w��96�9���9E4�9��9�99o�9z��9���9���9���9+��9hp�9��9���9�3�9ش�9�5�9P��9>�9��9x   x   B�9���9���9���9]��9��9�^�9���90�9٫�9@2�9���9+�9���9��9�N�9���9��9���9���9KM�9��9;��9�,�9ش�9^2�9}��9�2�9:��9�]�9x   x   L��9*��9���9��9���9G��9�N�9 ��9�)�9���9�5�9h��9�+�9���9z��9p,�9�X�9Fc�9rY�9�.�9%��9t��9�+�9���9�5�9v��9�&�97��9�Q�9���9x   x   �k�9�R�9�S�9�l�9���9��9�J�9���980�9Ӷ�9_3�9���9%�9�}�9���9� �9�9�9 �9���9'}�9��9@��9�4�9N��9�2�94��9I�9���9��9x   x   62�9y&�9�0�9{Z�99��9���9FP�9���9�?�9���9\4�9��9��9Fe�9C��9���9���9���9=��9)g�9�9��9j3�98��9>�9>��9�Q�9���9���9�Y�9x   x   �9�9T)�9�Z�9;��9���9�^�9���9�N�9��9;�9	��9��9E�9���9ߘ�9Y��9+�9/E�9� �9���9r;�9��9�P�9���9�]�9}��9��9�Y�9h)�9x   x   �D�9ZN�9sm�9M��9���9U+�9L��99��9:�9b��9���96:�9g�9&��9T��9���9���9���9��9@;�9q��9k��9�8�9c��9ׂ�9�*�9m��9��9�l�9QN�9x   x   UN�9<g�9��9��9���9hK�9��9��9�L�9��9���9l2�9�i�9���9���9+��9���94h�9-2�9���9���9�L�9p��9��9AK�99��9j��9&��9�f�9�M�9x   x   nm�9��9���9���9\'�9Gu�9���9��9�l�9���9B��91�9|Y�9�w�9�{�91x�9�Z�9b2�9���9���9kk�94�9���9{u�9�&�9b��9l��9H��9Tn�9_c�9x   x   6��9߸�9���93�9a�9���9���9�>�9���9X��9��9�.�9�N�9eZ�9nY�9�N�9W-�9\�97��9��9�A�9��9?��9�a�9��9���9t��9��9v��9���9x   x   ���9z��9Q'�9a�9Қ�9_��9O#�9�b�9P��9���9���9�(�9i>�9MA�9?�9G)�9���9���9���9�a�9"�9���9q��9b�9�%�9c��9M��9���9/��9���9x   x   ?+�9UK�9;u�9���9[��9r�9^Q�9w��9���9���9�
�9y(�9\2�9K2�9�'�9�
�9���9/��9���9NQ�9��9��9���9>v�96K�9[)�9V�9m
�9X�9S�9x   x   3��9���9���9���9K#�9]Q�9\�9ΰ�9���9���9��9@"�9�+�9�"�9}�9��9d��9���9@�9qQ�9!�9���9���9g��9z��9<f�9�V�9S�9gX�9�e�9x   x   ��9���9��9y>�9�b�9l��9ϰ�9^��9���9V�9��9
�9��9��9��9���9���9[��9!��9Ad�9�>�9��9���9N��9��9���9O��9Z��9��9G��9x   x   �9�9�L�9�l�9���9B��9���9���9���9��9q�9��9��9(�9C�9;�9[��9���9q��9:��9��9�j�9`L�9�:�9K'�9��9r�9~�9��9��9@&�9x   x   E��9���9���9F��9���9���9���9Q�9v�9�9j�9��9>�9��9��9"��9L��9u��94��9��9}��9.��9J��9Q��9�u�9�z�9 |�9�u�9���9z��9x   x   f��9���9/��9w�9���9z
�9��9��9��9d�9�9S�9��9��9��9�
�9���9��9���9c��9j��9���9/��9���9��9���9���9p��9���9���9x   x   :�9R2�91�9�.�9�(�9m(�97"�9�9��9��9Y�9��9��9k"�9�(�9�)�9`-�9-2�9�2�9R:�9]5�9iA�9�G�9�D�9�I�9eJ�9�F�9�F�9<@�9�5�9x   x   G�9�i�9dY�9�N�9\>�9T2�9�+�9��91�9>�9��9��9`*�93�9�<�9�O�9�Y�98h�9��9��9���9���9<��9±�9Y��9���9���9��9ї�9"��9x   x   	��9q��9�w�9]Z�9FA�9G2�9�"�9��9C�9��9��9s"�93�9B�9dZ�9�v�9P��9���9I��90��9���9E��9�9�9��9�90��96��9��9��9x   x   >��9���9�{�9eY�9?�9�'�9�9��9?�9��9��9�(�9�<�9_Z�92{�9[��9���9���9[�9r,�9�I�9�Z�9�o�9�q�9cn�9DZ�9J�9�.�9�9l��9x   x   ���9��9&x�9�N�9K)�9�
�9��9���9c��9.��9�
�9*�9�O�9�v�9[��9���9���9�0�93[�9���9���9n��9ü�9���9��9��9)��9RZ�9�0�9���9x   x   ���9���9�Z�9S-�9���9���9s��9���9���9^��9���9l-�9�Y�9d��9���9���9l<�9�u�9ß�9m��9���9;��92�9m��9���9���9���9�v�9=<�9&��9x   x   ���9)h�9f2�9\�9���9;��9��9l��9���9���9��9<2�9Hh�9���9���9�0�9�u�9u��9���9	�9�#�9�5�9I4�9U#�9i	�9���9ƫ�9�t�9d2�9���9x   x   ��9-2�9���9A��9���9���9Q�9>��9U��9M��9���9�2�9��9`��9f�9D[�9ʟ�9���9D�9�6�9�M�98[�91O�9i7�9Q�9���9���9�Y�9��9���9x   x   >;�9���9���9��9�a�9aQ�9�Q�9\d�9.��9��9{��9i:�97��9I��9�,�9ɂ�9y��9	�9�6�9�\�92m�9wm�9[�9~6�9�	�9���9Ղ�9�,�9���9?��9x   x   x��9���9wk�9�A�9$"�9��9!�9�>�9�j�9���9���95�9���9��9�I�9���9���9�#�9�M�92m�9q�9]m�9�O�9�#�9a��9ؚ�9�J�9���9���9�6�9x   x   u��9�L�9C�94��9���9!��9���9��9�L�9T��9���9�A�9���9e��9�Z�9���9M��9�5�9F[�9�m�9hm�9�Z�9k4�9s��9���9�X�9� �9���9\@�9���9x   x   �8�9}��9��9X��9���9���9��9���9�:�9o��9N��9�G�9b��91�9�o�9��9I�9Y4�9AO�9[�9�O�9i4�9V�9���9p�9,�9Ũ�92G�9���9'��9x   x   m��9'��9�u�9�a�9)b�9_v�9���9u��9u'�9���9���9�D�9��9E�9�q�9���9���9e#�9y7�9�6�9�#�9z��9���9�q�9��9���9{E�9m��9���9�'�9x   x   ނ�9NK�9�&�9��9�%�9YK�9���9)��9��9�u�97��9J�9~��9��9n�9���9���9	�9e�9�	�9g��9���9~p�9��9`��9?J�9���9�u�9S�9Y��9x   x   �*�9I��9x��9��9��9�)�9bf�9��9��9�z�9��9�J�9(��99�9dZ�9��9��9���9���9���9���9�X�96�9���9CJ�9���9�{�9��9n��9�d�9x   x   |��9x��9���9���9n��9v�9 W�9y��9��9L|�9���9�F�9���9R��9)J�9H��9Р�9׫�9ѡ�9��9�J�9� �9Ũ�9{E�9���9�{�9��9,��9Z�9��9x   x   ��92��9R��92��9���9�
�9%S�9~��9��9v�9���9�F�94��9X��9�.�9oZ�9�v�9�t�9 Z�9�,�9���9���92G�9h��9�u�9��9 ��9vP�9M	�9B��9x   x   �l�9�f�9bn�9���9L��9q�9�X�9��9�9���9	��9e@�9���95��9'�9�0�9Q<�9q2�9��9���9Ɩ�9_@�9���9���9Q�9k��9yZ�9E	�9:��9���9x   x   TN�9N�9kc�9���9���9l�9�e�9c��9g&�9���9��9�5�9H��9<��9���9���9:��9���9���9D��9�6�9���9&��9�'�9M��9�d�9��9<��9��9�d�9x   x   �t�9fz�9+��9��9F��9�)�9�k�9��9-�9�R�99��9���9|�9�-�9�L�9�Y�9�K�9�0�9��9���9���9�Q�95�9׻�9Gl�9J(�9:��9;��9��9Bz�9x   x   jz�9���9���9J��9|�9AA�9E��9��9��9p\�9\��9���9r�9|$�90�9�0�9�"�9��9���96��9&^�9�9#��9j��9�A�9@�9���9:��9M��9tz�9x   x    ��9���9���9c��9+�9
h�9���9)��9}1�9�p�9��9���9���9�	�9	�9�9���9j��9��9po�9h1�9���9���9]h�94*�9���9V��9&��9��9?��9x   x   ���9C��9_��9�!�9"S�9��9��9��9(F�9�x�9���9q��9{��9���9G��9��9Y��9���9�z�9�E�9��9���9��9iS�9�!�9���9r��9���9B��9��9x   x   =��9p�9+�9S�9x��9���9���9�-�9�[�9���9:��9,��9���9���9���9���9&��9���9[�9�,�9���9���9}��9�S�9�)�9�9��9@��9B��9���9x   x   �)�93A�9h�9��9���9���9|�99I�9�o�9���9���9���9���9���9���9i��9���9�n�9�J�9��9X��9���9Ð�9ih�9B�9�'�9�9��9g�9��9x   x   �k�91��9v��9��9���9{�9�D�9�j�9��9��9q��9U��9���9���9¹�98��9?��9<j�9�C�9w�9���9i��9��9���9�k�9�Z�9M�9-K�9�L�9�Y�9x   x   ��9��9��9��9�-�93I�9�j�9���9
��91��9C��9S��9Z��93��90��9��9 ��9�k�9I�9.�9��92��9���9ڻ�9���9t��9��9+��9u��9���9x   x   �9��9m1�9F�9�[�9�o�9��9��9Ӧ�9ݷ�99��9��9T��9���9��9���9$��9Gp�9iZ�9OF�9�0�9�9��9���9���9���9���9���9���9G��9x   x   ~R�9W\�9�p�9�x�9���9��9ޣ�9,��9��9���94��9l��9���9���9M��9��9��9��9Yy�9�p�9e]�9�R�9DH�9eA�9�>�9�5�9�7�9�?�9�@�9�H�9x   x   ��9H��9Ψ�9z��92��9���9p��9>��97��90��9U��9��9S��9L��9H��9���9%��99��9{��9��9B��9��9��9���9���9Z��9���9��9���9��9x   x   }��9u��9���9f��9"��9���9[��9M��9��9g��9��9���9��9i��9���9���9��9���9���9���9:��9���95��9���9���9���9��9��9���9���9x   x   b�9c�9���9l��9���9���9���9U��9T��9���9T��9��9���9���9S��9���9���9��9��9- �9�'�9�0�9]6�9�>�9/=�9�=�9�5�9�1�9#(�9V�9x   x   �-�9l$�9z	�9���9���9���9���9-��9Ŷ�9��9I��9e��9���9A��9���9c	�9�$�9�/�9@K�9�^�9�o�9�|�9�9���9Ň�9'��9G}�9�m�9L_�9YL�9x   x   �L�9 0�9��9F��9���9���9Ĺ�94��9��9X��9M��9���9[��9���9�	�9�/�9VK�9k�9���9"��9��9���9���9'��9��9���9��9���9a��9nk�9x   x   |Y�9�0�9�9 ��9���9a��9@��9 ��9���9���9���9���9���9k	�9�/�9�Z�9 ��9��9���9��9���9!�9��99�9<�93 �9���9��9��9Ѐ�9x   x   �K�9�"�9���9X��9+��9���9B��9��92��9���9.��9 ��9���9�$�9_K�9 ��9j��9���9���9��9y6�9[D�9D�9�D�9!6�9D�9R��9���9H��9���9x   x   �0�9��9f��9���9��9o�9Gj�9�k�9Sp�9���9K��9���9��9�/�9$k�9 ��9���9�	�9�3�9IM�99k�9�n�9�n�9k�9M�9�3�9��9z��9U��9�j�9x   x   ~�9���9��9�z�9![�9�J�9�C�9'I�9xZ�9ky�9���9��9��9LK�9��9���9���9�3�9sZ�9z�9���9���9���9�z�9Z�9�3�9��9y��9��9#J�9x   x   ���9>��9vo�9�E�9�,�9��9��9.�9`F�9�p�9��9��9F �9�^�94��9��9��9QM�9z�9Ք�9t��9���9��9�y�9�M�9��9��9���9�a�9��9x   x   ���9-^�9r1�9��9���9p��9���9��91�9�]�9_��9O��9(�9�o�9(��9���9�6�9Dk�9���9x��9(��9���9���9�j�9�6�9� �9@��9�l�9�&�9���9x   x   �Q�9�9���9���9���9���9~��9I��9.�9�R�9��9��9�0�9�|�9���94�9qD�9�n�9���9���9���9J��9�n�9�D�9��9���9�~�9�2�9���9��9x   x   D�9.��9���9%��9���9ݐ�9���9��9��9hH�9��9R��9}6�9݁�9���9��9D�9�n�9���9��9���9�n�9�D�9=�9���9���9R4�9���9d��9�I�9x   x   ��9x��9mh�9}S�9�S�9�h�9���9���9���9�A�9��9���9�>�9���9G��9T�9�D�9 k�9�z�9�y�9�j�9�D�9>�9��9j��9M@�9���9q��9r@�9���9x   x   Pl�9�A�9F*�9�!�9�)�9)B�9�k�9���9���9�>�9ё�9��9S=�9��9,��9Z�966�9M�9,Z�9�M�9�6�9��9���9k��9�<�9���9���9-?�9���9��9x   x   T(�9I�9���9���9�9(�9[�9���9���9�5�9��9���9>�9C��9���9I �9V�9�3�94�9��9� �9���9���9L@�9���9-��9�6�9���9Ԙ�9�Z�9x   x   E��9���9g��9���9#��9�95M�9<��9��9�7�9Ï�9%��9�5�9e}�9���9���9k��9��9#��9$��9N��9�~�9S4�9���9���9�6�9���9p��9,N�9��9x   x   G��9E��98��9׻�9R��9��9MK�9N��9���9�?�9/��9<��9�1�9n�9ڠ�9+��9���9���9���9���9�l�9�2�9���9p��9*?�9���9r��9?I�9��9g��9x   x   ��9P��9���9P��9Q��9��9�L�9���9���9�@�9ܕ�9���9?(�9d_�9}��9��9Y��9d��9��9�a�9�&�9���9`��9m@�9���9Θ�9,N�9��9B��9���9x   x   Dz�9wz�9N��9��9���9��9�Y�9ۧ�9_��9�H�9;��9���9r�9pL�9�k�9��9���9�j�9+J�9��9���9'��9�I�9���9��9�Z�9��9`��9���9���9x   x   W{�9N��9���9j��9���9I�9�V�9���9��9B�9�F�9P{�9���9r��9���9h��9��9y��9E��9�z�9CF�9��9���9f��9�U�9Q�9;��9ƺ�9���9��9x   x   O��9���9��9���9���9�3�9	o�9��9���9��9TK�9<x�9j��9���9���9���9���9Y��9!x�9�L�9P�9���9ۜ�9�n�95�9J��9���9���9��9��9x   x   ���9��9c��9���9��95N�9Ђ�9���9���9w%�9=Q�9�s�9���9���9��9���9���9�t�9�P�9�#�9���9l��9���9N�9��9��9���9=��9��9��9x   x   h��9���9���9.�9B�9kl�9\��9��9o��9X.�94P�98v�9ш�91��9��9���9�u�98O�9!0�9���9
��9��9�l�9-B�9��9���9 ��9���9��9��9x   x   ���9���9��9B�9�k�9*��9���9Q��9��9?<�9�[�9zs�9/|�9���9	~�9�s�9s\�9"<�9��9���9$��9_��9qk�9YB�9��9@��9���9Z��9��9/��9x   x   ;�9{3�9*N�9dl�9(��9N��9���9#�9*�9�I�9�Z�9xl�9r|�9|�9�j�9hZ�9�I�9�)�9��9���9ִ�9���9Il�9iM�9�4�9��9I�9��9*�9��9x   x   �V�9�n�9ł�9Z��9���9���9��9p�9n;�9[Q�9�\�9!m�9�q�9\m�9�^�9mP�9<�9Y�9��9��9O��9��9��9n�9�U�9nF�9�<�9�=�9�;�9E�9x   x   ��9u��9���9��9I��9 �9q�9�7�9�O�9V]�9�f�9qf�99f�9f�9�\�9�O�9H7�9��9%�9���9&��9���9���9T��9��9�u�9t�9Lu�9�w�9���9x   x   ��9���9���9b��9��9
*�9i;�9�O�9GX�9@^�9mg�9�f�9;h�9�]�9�Y�9$O�9�;�9�*�9��9��9G��9I��9*��9���9c��9��9ʲ�9c��9*��9}��9x   x   /�9��9b%�9I.�93<�9�I�9]Q�9W]�9<^�9�b�9<h�9Vg�9�b�95^�9k\�97R�9�G�93<�9C0�9�#�9?�9&�9#�9� �9|��9��9q��9���9���9b�9x   x   �F�9EK�9.Q�9/P�9�[�9�Z�9�\�9�f�9jg�9Bh�9 k�9<h�9[g�9�f�9�\�9�[�9�]�9�M�9jQ�9ML�9�E�9�G�9@�9kA�9:E�9^G�9�B�9B�9a@�9RG�9x   x   6{�9%x�9�s�9,v�9ps�9kl�9m�9rf�9�f�9[g�9?h�9Gf�9�f�9tn�9*j�9rq�9*w�9Pt�9�w�9�{�9���9-��9+��9	��9	��9��9υ�9g��9���9+��9x   x   ��9[��9���9ˈ�91|�9k|�9�q�9:f�99h�9�b�9[g�9�f�9�o�9}�9��9!��9i��9���9��9���9���9¿�9X��9���9[��9���9���9K��9E��9W��9x   x   [��9���9{��9!��9��9{|�9Zm�9f�9�]�9=^�9�f�9|n�9}�9-��9א�9Ρ�9���9L��9���9h��9���9��9��9	�9�9��9��9���9���9.��9x   x   ���9���9��9��9~�9�j�9�^�9�\�9�Y�9k\�9�\�96j�9��9ݐ�9%��9���9���9��9�
�9h$�9�/�9yA�9�E�9J�9�F�9g@�9�/�9S%�9��9��9x   x   X��9���9���9}��9�s�9jZ�9sP�9�O�9-O�97R�9�[�9zq�9!��9ӡ�9���9Z��9{�9R�9�?�9sT�9*c�9�y�9>}�9�|�9�y�9�c�9�S�9@�9��9�9x   x   ���9��9���9�u�9u\�9�I�9 <�9X7�9�;�9�G�9�]�99w�9o��9���9���9t�9�(�9�M�9Xn�9@��9r��9��9~��9���9^��9`��9an�9�M�9D'�9��9x   x   w��9[��9�t�9:O�9&<�9�)�9g�9��9�*�9C<�9�M�9bt�9���9]��90��9X�9�M�9�r�9��9s��9���9A��94��9/��9Ʈ�9O��9�r�9�M�9��9���9x   x   A��9x�9�P�9&0�9��9��9��92�9�9Y0�9yQ�9�w�9)��9���9�
�9�?�9`n�9���9���9��9���9���9U��9���9���9���9�n�9�@�9 	�94��9x   x   ~z�9�L�9�#�9 �9 ��9���9��9���9-��9�#�9`L�9�{�9���9}��9t$�9�T�9N��9w��9"��9h��96��9��9���9���9��9A��90S�96%�9���91��9x   x   JF�9V�9���9��93��9��9a��97��9_��9N�9�E�9���9���9��9�/�97c�9}��9���9���9@��9}��9K��9���9O��9��9�d�9�/�9���9���9���9x   x   ��9���9~��9���9o��9͔�9��9���9g��9A�9�G�9G��9տ�9��9�A�9�y�9���9J��9���9��9K��9]��9���9���9�x�9*@�9��9c��9^��9�G�9x   x   ���9���9��9�l�9�k�9]l�9%��9�9F��9D�9;@�9E��9u��9��9�E�9O}�9���9B��9`��9���9���9���9 ��9X}�9�G�9��9���9���9�?�9i�9x   x   i��9�n�9$N�99B�9iB�9}M�9%n�9i��9���9� �9�A�9��9���9 �9�J�9�|�9���9<��9���9���9W��9���9P}�9�I�9d�9���98��9+B�9���9���9x   x   �U�95�9��9��9��9�4�9�U�9��9���9���9VE�9"��9y��9�9	G�9�y�9r��9֮�9���9��9��9�x�9�G�9b�9d��9��9dC�9v��9���9V��9x   x   \�9U��9)��9���9Y��9��9�F�9�u�9��9;��9xG�9���9 ��9��9}@�9�c�9t��9_��9���9J��9�d�9+@�9��9���9��9�H�9:��9���9sv�9�G�9x   x   @��9���9���9��9���9d�9�<�90t�9��9���9C�9��9���9��9�/�9�S�9rn�9�r�9�n�9:S�9�/�9��9���9>��9eC�97��9���9qu�9�;�9Z�9x   x   Һ�9���9L��9��9l��9��9�=�9du�9~��9���9$B�9���9c��9���9g%�9@�9�M�9�M�9�@�9<%�9���9g��9���93B�9u��9���9uu�9=�9��9���9x   x   �9��9��9��9&��9<�9<�9�w�9B��9���9}@�9���9]��9���9��9��9R'�9��9	�9���9���9[��9�?�9���9���9nv�9�;�9��9���9o��9x   x   $��9���9��9���9E��9��9(E�9ւ�9���9z�9iG�9B��9j��9=��9(��9�9��9���9;��9;��9���9�G�9b�9���9W��9�G�9U�9���9r��9���9x   x    ��9A��9���9M��9���9��9�0�9�f�9���9g��9 ��9((�91H�9b�9Wq�9Fy�9#p�9�a�9:I�9�&�9���9���95��9�h�9N/�9� �9��9���96��9��9x   x   A��9��9{��9���9I��9�9�C�9 x�9���9���9E��9v#�9�=�9�M�9h_�9�_�9�N�9�=�9�"�9r��9��9���9�u�9]C�9G�9n��9%��9��9c��9��9x   x   ���9x��9���9���9��9-(�9�X�9{��9��9x��9���9K�9<4�9TB�9xH�9�A�9�3�9��9# �90��9��9+��9�Y�9?'�9��9d��9@��9���9S��9���9x   x   E��9���9���9���9S �9{F�9�m�9�9���9���9��9�9/�9�4�9�4�9�/�9M�9��9���9b��9f��9�l�9�F�9� �98��9���9x��9´�9U��9I��9x   x   ���9E��9��9P �9�B�9Nc�97��9S��9��9��9r��9T�9"�9P!�9�!�9�9j��9��9���9^��9���9�b�9�B�9w �9 �9O��9@��9���9��9��9x   x   ��9�9)(�9yF�9Ic�9/��9!��9p��94��9���9R�9/�9��9��9'�9��9O��9v��9���9��9���9Vd�9�E�9�&�9C�9��9���94��9��9���9x   x   u0�9�C�9�X�9�m�94��9 ��9c��9F��9t��9���91�9��9d�9[�9��9:��9;��9y��9���9��9Ɇ�9�l�9�Z�9C�9�/�9�#�9��9l�9M�9$#�9x   x   �f�9�w�9j��9���9L��9m��9C��9Z��9:��9��9%�9(�9l�94�9i�9���9/��9?��9P��9
��9ǚ�9#��95w�9lg�9jW�9�Q�9(H�9[H�9NR�9�V�9x   x   n��9���9��9���9��93��9r��99��93�9Y�9s�9�9��9��9��9���9���9��9���9��9<��9���9���9���9`��9x��9#��9���9��9���9x   x   W��9}��9j��9���9���9���9���9��9U�9��9^�9��9n�9o�9J�9<��9t��9���9���9+��9c��9���9���9���9���9��9ܹ�9b��9N��9��9x   x   ��95��9���9��9f��9Q�9,�9(�9r�9^�9�9v�9h�9��9'�9��9� �9"�9X �9P��9=��9!��9E��9��9?��9���9X��9���9���91��9x   x   (�9l#�9B�9��9L�9.�9��9,�9�9��9x�9��9��9��9W�9�9��9��9"�9�&�9�"�9�'�9�.�9
)�9-�9�-�9�)�9�.�9'�9�"�9x   x   $H�9�=�904�9/�9"�9��9d�9p�9��9m�9j�9��9��9X�9�$�9=.�9A3�9>�9VI�9�P�9�V�9�[�9�a�9�e�9ue�9�e�9�`�9,\�9iW�9TO�9x   x   b�9�M�9JB�9�4�9I!�9��9T�9:�9��9o�9��9��9[�9��9j4�9C�9�M�9�a�9gp�9��9ǋ�9ʍ�9���9)��9P��9x��9Ɏ�9���9l��9�q�9x   x   Qq�9Y_�9rH�9�4�9�!�9%�9��9j�9��9P�9*�9S�9�$�9i4�9!H�9?_�9q�9���9)��9"��9���9��9���9���9���9���9Ķ�9���9ē�9Q��9x   x   >y�9�_�9�A�9�/�9 �9��99��9���9���9B��9��9�9C.�9%C�9F_�9wy�9ڎ�9ߧ�9��9���9f��9���9���9x��9P��9���9U��9���9���9���9x   x   !p�9�N�9�3�9L�9k��9S��9>��9/��9���9}��9� �9��9J3�9�M�9q�9ڎ�9���9g��9v��97�9��9��9t�9��9v�9�9���9���9]��9���9x   x   �a�9�=�9��9��9���9��9���9E��9��9���9+�9��9>�9�a�9Ã�9��9m��98��9��9�!�9-*�9(1�9U2�9�*�9�!�9t�9���9���94��9I��9x   x   :I�9�"�9- �9���9���9���9���9]��9���9���9f �9"�9fI�9pp�9,��9���9x��9��9�"�9�6�9C�9>H�9�A�97�9�!�9��9<��9��9���9�p�9x   x   �&�9p��94��9j��9i��9���9��9��9��9=��9a��9�&�9�P�9 ��9(��9���9;�9�!�9�6�9�L�9�V�9RW�9�L�9�6�9�"�9��9���95��9��9cP�9x   x   ���9��9���9i��9��9���9Ն�9Ӛ�9I��9p��9R��9#�9�V�9ڋ�9���9v��9��93*�9C�9�V�9�W�9�V�9�B�9�)�9�9��9F��9 ��9#W�9K#�9x   x   ���9���92��9�l�9�b�9fd�9m�98��9���9���94��9�'�9�[�9ݍ�9��9���9��941�9BH�9TW�9�V�9YH�9	2�9d�9*��9;��9k��9�\�9 '�9���9x   x   6��9�u�9�Y�9�F�9�B�9F�9[�9Ew�9��9���9U��9�.�9�a�9���9���9���9��9c2�9�A�9M�9�B�92�95�9��9���9���9�`�9y.�9f��9���9x   x   �h�9fC�9J'�9� �9� �9'�9-C�9�g�9�9��94��9$)�9�e�9<��9���9���9�9�*�97�9�6�9�)�9g�9��9U��9Ԙ�99e�9T*�9��9��9���9x   x   R/�9J�9��9B��9/�9P�9�/�9W�9t��9ҵ�9W��9-�9�e�9h��9��9b��9��9�!�9�!�9#�9�91��9���9֘�9f�9c-�9;��9F��9ރ�9V�9x   x   � �9x��9t��9���9]��9��9�#�9�Q�9���9��9���9�-�9�e�9���9���9	��9�9�9��9��9��9A��9���9:e�9f-�9���9i��9��9-R�9Z%�9x   x   ��9.��9P��9���9O��9���9��9AH�9:��9��9n��9�)�9�`�9ݎ�9׶�9l��9��9���9G��9���9I��9n��9�`�9L*�99��9m��9���9�H�9��9O��9x   x   ���9��9���9ϴ�9���99��9��9qH�9��9x��9��9�.�9A\�9���9���9ȿ�9���9���9���9;��9"��9�\�9y.�9���9E��9��9�H�9��9��9���9x   x   :��9n��9Y��9]��9-��9��9c�9^R�9"��9c��9���9.'�9W�9���9ғ�9Ԩ�9i��9>��9���9��9*W�9
'�9g��9��9݃�9-R�9��9 ��9��9Ԭ�9x   x   ��9��9���9M��9"��9���99#�9�V�9���9 ��9D��9#�9bO�9�q�9\��9���9���9S��9�p�9^P�9N#�9���9���9}��9 V�9W%�9G��9���9Ь�9��9x   x   ���9�|�9��9٤�9ӿ�9��9�9L-�9�W�9M�9o��9���9>��9���9�
�9��94
�90��9���96��9M��9~��9�W�9-/�9��9���9��9���9a��9U|�9x   x   �|�9E��9͙�9��9 ��9���9g�9;>�9�b�9���9���9k��9���9m��9��9��9���9 ��9���9���9!��9Cc�9�;�9�9���9���9���9	��9���9�z�9x   x   ��9Ι�9"��9G��9z��9|�9M'�9$I�9�o�96��9���9��9���9���9{��9Y��9���9���9̭�9��9�o�9 K�9�(�9��9���9(��9¬�9���9g��9���9x   x   Ϥ�9��9D��9K��9���9��9�7�9�\�9}�9��9Ķ�9���9V��9A��9���9;��9���9���93��9H�9Z�9S6�9D �9T��9���9���9[��9ʣ�9���9���9x   x   ʿ�9���9r��9���9�9t3�9�N�9Lr�9��9��9���9���9���9���9���9ֿ�9 ��9��9��9yr�9�Q�9j2�9��9���9��9=��9Y��9���9.��9��9x   x   ��9���9~�9��9k3�9JQ�9ae�9��9��9q��9^��9C��9��9���9(��9t��9٫�9���9a�9�c�9`P�9�4�9��9��9���9��9���9���9���9���9x   x   v�9\�9J'�9�7�9�N�9de�9�v�9��9Q��9~��9��9��9���9���9Q��9��9���9,��9�x�9�e�9�N�9�6�9s)�9��9(�9���9���9���9^��9��9x   x   >-�94>�9I�9�\�9Hr�9��9��9u��9~��9��9y��9���9���9`��9)��9Э�9���9���9y�9�r�9�\�9_H�9:=�9�,�9P&�9� �9'�9s�9��9&�9x   x   �W�9�b�9�o�9�|�9��9��9O��9���9��9O��9T��9|��9ķ�9���9j��9H��9���9���9���9�|�9�q�9�b�9TY�9dN�9jJ�9	G�99D�9\G�9FK�9O�9x   x   >�9���9.��9��9��9n��9w��9���9O��9.��9J��9>��9��9%��9	��9ʮ�9���9I��9��9J��9q��9�~�9�|�9"{�9h|�9�s�9�s�9]|�9�y�9�}�9x   x   a��9���9���9���9���9Z��9��9x��9V��9K��9w��9{��93��9���9���9���9	��9���9N��9���9^��9��9���9Z��9J��9~��9a��9��9���9���9x   x   ���9]��9���9���9���9C��9��9���9y��9<��9u��9��9���9���9��9��9���9���9p��96��9��9��9_��9���9x��9���9���9���9��9���9x   x   .��9���9���9P��9���9��9���9���9Ƿ�9"��96��9���9���9���9G��9���9��9���9���9���9���9f��9A��9��9��9��9Q��9���9��9	��9x   x   ���9d��9���9C��9���9���9���9`��9���9'��9���9��9���9���9i��9���9P��9���9
�9��9�9v$�9(�9 '�9�&�9I*�9�$�9��9��9`�9x   x   �
�9��9s��9���9���9*��9S��92��9o��9��9���9��9Q��9e��9���9\��9��9J�9p/�9�2�9�F�9�O�9�T�9IV�9�S�9*N�9�G�9 3�9�.�9��9x   x   t�9 ��9N��9?��9ֿ�9t��9��9ӭ�9K��9Ԯ�9���9"��9���9���9U��9��9�&�9�A�9�N�9�^�9�l�9�r�9Y{�9�{�91t�9�l�9�]�9�O�9�A�9�&�9x   x   3
�9���9���9���9��9٫�9���9���9 ��9���9��9���9��9Z��9��9�&�9�9�9Q�9mi�9�v�9m��9���9���9ߔ�9��9'v�9Ji�9�O�9J:�9!'�9x   x   ,��9���9���9���9��9���93��9��9���9V��9ϴ�9���9���9���9Q�9�A�9Q�9x�9��9��9���9Ѭ�9���9���9���9���9mx�9�Q�9r@�9��9x   x   ���9���9ɭ�90��9��9b�9�x�9}�9���9���9Z��9��9���9
�9w/�9�N�9si�9��9���9��9��9���9o��9u��9��9։�9xi�9�N�9�/�9��9x   x   /��9���9��9M�9}r�9�c�9�e�9�r�9�|�9U��9��9<��9���9��9�2�9�^�9�v�9��9��9#��9,��9F��9S��9>��96��9Zw�9~]�9$4�9>�9���9x   x   L��9'��9�o�9Z�9�Q�9jP�9�N�9�\�9�q�9���9n��9���9���9�9�F�9�l�9x��9���9��9.��9��9#��9���9��9ۅ�9�m�9^F�9��9"��9^��9x   x   ���9Mc�9$K�9\6�9u2�9�4�97�9kH�9�b�9�~�9��95��9{��9�$�9�O�9�r�9���9ܬ�9���9F��9%��9��9j��9���9Ns�9�O�9m#�96��9.��9Y��9x   x   �W�9�;�9�(�9K �9��9��9z)�9I=�9dY�9�|�9���9k��9N��9�(�9�T�9b{�9 ��9í�9u��9P��9���9n��9ޒ�9�{�9WS�9o*�9��9���9ʦ�9|�9x   x   -/�9 �9��9c��9���9��9��9�,�9vN�97{�9h��9���9��9'�9RV�9�{�9��9���9|��9G��9
��9���9�{�9�V�91'�9��92��9���9�z�9*O�9x   x   ��9���9���9���9��9���98�9\&�9J�9x|�9Z��9���9��9'�9�S�9?t�9���9˒�9��9?��9���9Os�9US�90'�9��9���9���9*|�97K�9�$�9x   x   ���9���91��9���9N��9.��9���9� �9G�9�s�9���9���9
�9Y*�9<N�9�l�9-v�9��9؉�9[w�9�m�9�O�9j*�9��9���9��9�t�9G�9� �93��9x   x   ���9���9̬�9d��9f��9���9���92�9OD�9	t�9s��9���9b��9�$�9�G�9^�9Ti�9x�9i�9�]�9fF�9q#�9"��96��9���9�t�9JC�92�9��9N��9x   x   ���9��9��9գ�9���9���9���9|�9pG�9o|�9,��9���9���9��93�9�O�9�O�9�Q�9�N�9(4�9��92��9���9���9*|�9G�9.�9���9/��9���9x   x   f��9ȃ�9r��9���9@��9��9o��9��9YK�9�y�9Ȥ�9 ��9��9��9�.�9�A�9P:�9|@�9�/�9A�9#��9&��9Ǧ�9�z�99K�9� �9��94��9���9W��9x   x   M|�9�z�9���9���9��9���9��9&�9O�9�}�9���9���9��9s�9��9�&�9+'�9��9��9���9a��9S��9|�9*O�9�$�9-��9Q��9���9T��9V��9x   x    f�9�i�9�r�9��9��9��9���9��9��9F?�9C[�9Dy�94��9H��9���93��9���9"��9H��9�w�9b\�9�@�9��9 ��9B��9j��9���90��9+q�9si�9x   x   �i�9�o�9�|�9��9���9���9���9A�9�&�9�D�9s^�9'z�9U��9=��9=��9ܞ�9���9��9�y�9�^�9�B�9�&�9|�9���9<��91��9	��9g}�9�p�9ah�9x   x   �r�9�|�9`��9h��9���9��9��9��9#+�9�M�9Vb�9v�9��9���9���9N��91��9u�9c�9^N�9e+�94�9���9���9���9`��9$��9�{�9cs�94s�9x   x   ��9��9f��9���9y��9���9��9��9�2�9�P�9^�9
v�9�~�9��9r��9W�9lw�9J^�9�N�9
4�9b�9��9���90��9��9���9��9�~�9��9O�9x   x   ܚ�9���9���9v��9N��97��9��9(+�9|C�9�V�9.d�9�u�9�x�9�s�9�v�9u�9�b�9{X�9�B�9Q+�9��9Q��9���9���9+��9-��9Ú�9���9��9Ò�9x   x   ��9���9��9���91��9f	�9!�9B;�9�J�9HW�9	`�9�n�9Cw�9�v�9�p�9a�9�U�9�J�9 ;�91 �9��9o��9M��9E��9���9)��9K��9��9���9���9x   x   ���9���9��9��9��9!�938�9D�9�Q�9�\�9�g�9�o�9jn�9(p�9�d�9�^�9(Q�9JD�99�9!�9��9��9X��9C��9d��9{��9J��9���9l��9M��9x   x   ��98�9��9��9%+�9C;�9D�9�O�9�[�9�c�9n�9�k�9Hk�9uo�9�c�9e[�9{P�9�B�9];�9h+�9)�9�9�9���9`��9���9���9��9��9���9x   x   ��9�&�9+�9�2�9uC�9�J�9�Q�9�[�9`�9g�9�j�9�m�9�i�9�h�9(_�9�[�9"R�9K�9�B�9e2�9�,�93&�9�9��9��9N	�9s�9�
�9�9��9x   x   9?�9�D�9�M�9�P�9�V�9CW�9�\�9�c�9g�9kl�9�m�9Yp�9�j�9Mf�9�e�9�[�9W�9}V�9�Q�91L�9�C�9�?�9�:�9�4�9�/�9�2�9J1�9�/�9�4�9	;�9x   x   >[�9n^�9Rb�9
^�9'd�9�_�9�g�9n�9�j�9�m�96e�9*n�9m�9`m�9�f�9�`�9�c�9]�9�b�9'`�9s[�91[�9�V�9�U�9X�9I\�9-X�9'V�9�U�9 \�9x   x   5y�9z�9v�9v�9�u�9�n�9�o�9�k�9�m�9[p�9&n�9�l�9�j�9Dp�9�o�9u�9�w�9�u�9�x�9�w�9�{�9�z�9��9~�9dy�9�z�9�}�9��9�z�9�z�9x   x   ,��9M��9��9�~�9�x�9Aw�9hn�9Kk�9�i�9�j�9m�9�j�9�o�9v�9Yx�9~�9ă�9l��9{��9���9���9��9���9���9���9���9ģ�9��9*��9<��9x   x   ?��94��9}��9w�9�s�9�v�9(p�9so�9�h�9Nf�9am�9Hp�9v�9Yt�9���9`��9I��9���9���9մ�9���9+��9��9���9���9���9���9μ�9}��9��9x   x   ���9?��9z��9h��9�v�9�p�9�d�9�c�9)_�9�e�9�f�9�o�9Sx�9���9���9k��9H��9���9W��9x��9���9���9���9���9?��9	��9p��9/��9���9���9x   x   ,��9ݞ�9N��9S�9u�9a�9�^�9d[�9�[�9�[�9�`�9u�9~�9g��9h��9?��9���9I��9$��9���9��9���9b��9���9��9X��9���9���9;��9���9x   x   ��9���9-��9jw�9�b�9�U�91Q�9�P�9'R�9�W�9�c�9�w�9ƃ�9Q��9H��9���9���9���9Y��96�99�9Z�9�9��9��9�
�95��9K��9���9���9x   x   ��9���9u�9P^�9~X�9�J�9OD�9�B�9K�9�V�9
]�9	v�9s��9���9���9L��9���9J �9�9&!�9G(�9-�9.�92(�9�!�9��9 �9��9	��9I��9x   x   A��9�y�9c�9�N�9C�9;�9#9�9b;�9�B�9�Q�9�b�9y�9��9���9^��9'��9\��9�96%�9�1�9�7�9�=�97�92�9?$�9)�9���9��9���9w��9x   x   �w�9�^�9aN�94�9U+�97 �9!�9q+�9s2�9=L�9/`�9�w�9˖�9۴�9���9���9:�9#!�9�1�9g9�9�D�9�D�9�9�9�1�9�"�9��9]��9���9���9���9x   x   e\�9�B�9g+�9i�9��9��9��91�9�,�9�C�9~[�9�{�9���9���9���9��9>�9J(�9�7�9�D�9YK�9�D�9J7�9�'�9!�9���9���98��9���9O{�9x   x   �@�9�&�96�9��9]��9|��9�9"�9=&�9�?�9;[�9�z�9��96��9���9���9f�9-�9�=�9�D�9�D�9�=�9�-�9��9���9���9���9��9�z�9�Z�9x   x   ��9��9���9���9���9[��9i��9/�9-�9�:�9�V�9��9���9��9���9q��9�9.�97�9�9�9K7�9�-�9>�9���9���9?��9��9G�9�W�9�9�9x   x   ��9���9���95��9��9S��9O��9���9��9�4�9�U�9~�9��9���9���9���9��95(�92�9�1�9�'�9��9���9&��9���9���9�}�9�T�9�5�9T�9x   x   H��9B��9���9��92��9���9q��9s��9��9�/�91X�9oy�9���9���9M��9%��9��9�!�9A$�9�"�9&�9���9���9���95��9�z�9�Y�9�.�9m�9\��9x   x   n��96��9h��9���96��9:��9���9���9]	�9�2�9V\�9�z�9à�9���9��9d��9�
�9��9/�9��9���9���9A��9��9�z�9qY�9�2�9�	�9���9���9x   x   ���9��9*��9��9̚�9X��9W��9���9��9U1�9=X�9�}�9ӣ�9���9{��9���9<��9 �9���9b��9���9���9��9�}�9�Y�9�2�98�9b��9'��95��9x   x   6��9o}�9�{�9�~�9��9��9���9-��9�
�9�/�97V�9��9$��9ۼ�9>��9���9T��9 ��9��9���9:��9��9C�9�T�9�.�9�	�9e��9���9E��9��9x   x   /q�9�p�9fs�9��9#��9���9r��9'��9�95�9�U�9�z�9;��9���9���9D��9���9��9���9���9�9�z�9�W�9�5�9f�9���9"��9=��9y��9��9x   x   |i�9ih�9:s�9V�9ǒ�9ǭ�9V��9���9��9;�9\�9�z�9K��9��9��9���9���9N��9{��9���9N{�9�Z�9�9�9T�9W��9���9/��9��9��9Ht�9x   x   ?�9dI�9�R�9Fa�9�u�9r��9��9Ž�9���9���9R�9f*�9:7�9�I�9$S�9YU�9#S�9jG�9�6�9k)�9_�9���9K��9��9���9��9au�9ka�9�P�9@I�9x   x   bI�9�Q�9
W�9�k�9v�9-��9��9���9c��9f��9��9$�9>2�9:�9�E�9�D�9�;�93�9�$�9��9,��9���9���9Y��9Q��9&�9�k�9�W�9NS�9HI�9x   x   �R�9W�9�_�9 v�9���9��9���9c��9H��9f��9��9%'�9�1�9�4�9H>�9s4�9�0�9&�9�9���9��9I��9��9���9���9�v�9�^�9V�9�Q�9aL�9x   x   Ca�9�k�9�u�9Ǉ�9:��9`��9Q��9���9k��9%�9��9�!�9�+�981�9r2�9�+�9m#�9��9��9���9(��9���9���9���9��9bv�9�m�9^a�9�X�9X�9x   x   �u�9u�9���9?��9���9��9���9���9��9��96�9�!�9�'�9�,�9�&�9g!�9�9��9���9���9=��9��9��9���9��9�}�9�t�9;m�9�l�9�l�9x   x   j��9#��9��9d��9 ��9���9/��9
��9� �9X�9��9� �9�#�9�#�9�!�9��9k�9a �96��9���9���9���9h��9���9)��9���9u��9�{�9_}�9��9x   x   ޜ�9��9���9L��9���9*��9$��9� �9�9_�9e�9��9��92�9o�9��96�99�9&��9e��9_��9��9v��9>��9Ŝ�9W��9͚�9 ��9���9��9x   x   ���9���9^��9���9���9	��9� �9G�9��9B�9��9��9`�9��9��92�9Y	�9�9~��9���9��9���9T��9о�9`��9 ��9���9���9n��9*��9x   x   ���9]��9H��9g��9��9~ �9�9��96�9)�9@�9| �9�9��9��9��9��9� �9x��9���9���9���9���9��9���9E��9��9Y��9��9��9x   x   ���9]��9Z��9�9��9V�9`�9?�9+�9O�9w�9��9��9��9I�9��9G�9i�9A�9��9I��9���98��9C��9B��9���9��9���9���9���9x   x   I�9��9��9��97�9��9a�9��9=�9q�9��9z�9�9��9��9s�9��9v�9��9U�9�9�
�9D�9_�9j	�9:�9�	�9�9�9��9x   x   ^*�9$�9'�9�!�9�!�9� �9��9��9v �9��9}�9 �9��95�9� �9�!�9I#�9I&�9Q$�9�*�9�*�9M(�9/�9v-�9�.�9�/�9�,�9�/�9)�9	*�9x   x   17�922�9�1�9�+�9�'�9�#�9��9]�9�9��9�9��9��9O#�9(�9�*�9�0�9�2�9�5�9�=�9VB�9�A�9yE�9�I�9�K�9I�95F�9.A�9B�9�=�9x   x   I�9�9�9�4�921�9�,�9�#�92�9��9��9��9��93�9P#�9�,�9�1�9�5�9K:�9�I�9�M�9�W�9T]�9^a�9^c�9�c�9�c�9�c�9�`�9x]�9vX�9M�9x   x   S�9�E�9C>�9n2�9�&�9�!�9j�9��9��9N�9��9� �9(�9�1�9�=�9LE�92R�9;]�9�e�97s�9st�9~��9D��9�}�9���9��9�u�9Xr�9�e�9�\�9x   x   PU�9�D�9w4�9�+�9j!�9��9��91�9��9��9r�9�!�9 +�9�5�9SE�9SV�9^c�9�m�9hz�9m��9��9L��9ƛ�9���9ߚ�9���9��9nz�9mn�9Ec�9x   x   S�9�;�9�0�9o#�9�9t�98�9Z	�9��9Q�9��9S#�9�0�9L:�94R�9]c�9�x�9���9��9���9��9G��9k��9c��9��9A��9���96��9�x�9hc�9x   x   jG�93�9&�9��9��9a �9<�9�9 �9k�9x�9T&�9�2�9�I�9>]�9�m�9���9L��9���9��9���9q��9��9ӳ�9��9���96��9>��9�m�9�]�9x   x   �6�9�$�9�9��9���9B��9.��9���9~��9K�9��9W$�9�5�9�M�9�e�9iz�9��9���9S��9��9��9���9���9��9���9M��9K��9�z�9Le�9�N�9x   x   l)�9��9���9���9���9���9m��9���9���9��9^�9�*�9�=�9�W�99s�9q��9���9��9��9k��9���9���9���9���9Y��9��9ւ�9|s�9dV�92>�9x   x   a�90��9&��9,��9F��9���9j��9!��9���9U��9)�9�*�9`B�9`]�9zt�9���9��9���9��9���9���9���9Z��9���9b��9���9Qt�9_�9xB�9&*�9x   x   ���9���9O��9���9
��9���9��9��9���9���9�
�9O(�9�A�9ja�9���9P��9L��9t��9���9���9���9i��9���9���9l��9<��9�_�9�@�9%)�9t
�9x   x   N��9���9��9ˮ�9���9o��9|��9Z��9���9E��9Q�9/�9�E�9ic�9N��9˛�9p��9��9���9���9Z��9���9
��9+��9�~�9�d�9kG�9^/�9\�9O��9x   x   ��9]��9���9���9���9���9G��9޾�9��9N��9j�9�-�9�I�9 d�9�}�9���9n��9ڳ�9���9���9���9���9+��9�~�9�c�9�G�9�,�9	�9���9���9x   x   ���9U��9���9��9��93��9Μ�9o��9��9O��9u	�9�.�9�K�9�c�9���9��9$��9��9Ű�9\��9d��9p��9�~�9�c�9M�9�/�95�9B��9��9���9x   x   ���9+�9�v�9mv�9�}�9��9[��9&��9K��9���9K�9�/�9 I�9�c�9��9���9K��9���9X��9��9���9B��9�d�9�G�9�/�9/�9O��9���9ʲ�9���9x   x   cu�9�k�9�^�9�m�9�t�9���9ٚ�9���9��9)��9�	�9�,�9CF�9a�9�u�9��9��99��9T��9ڂ�9Rt�9�_�9nG�9�,�98�9S��9���9w��9��9 ��9x   x   pa�9�W�9)V�9ia�9Dm�9�{�9-��9���9b��9���9�9�/�9;A�9]�9\r�9sz�9@��9>��9�z�9�s�9_�9�@�9]/�9�9F��9���9y��9ѕ�9}�9�l�9x   x   �P�9HS�9�Q�9�X�9�l�9d}�9���9x��9��9���9�9$)�9B�9~X�9�e�9vn�9�x�9�m�9Oe�9`V�9xB�9+)�9\�9���9��9̲�9��9}�9pk�9)Y�9x   x   FI�9MI�9`L�9&X�9�l�9���9%��96��9��9���9��9*�9�=�9M�9�\�9Gc�9lc�9�]�9�N�9->�9$*�9w
�9M��9���9���9���9���9�l�9(Y�9;M�9x   x   �$�9"�9J)�9�7�9P>�9�Y�9,m�9#��9;��9��9s��9���9���9���9m��9���93��9���9���9z��9���9���9ޛ�9˅�9jm�9�Z�9#=�9m7�9f(�9	"�9x   x   "�9V!�9 2�9&7�9�K�9�a�9�p�9���9���9ص�9y��94��9h��9c��9+��9���9��96��9��9P��9M��9:��9���9q�9E`�9%L�9�7�9�2�9�!�9$"�9x   x   G)�9�1�9�<�9-H�9.X�9l�9}�9��9���9ַ�9���9���95��9i��9��9���9}��9��9J��9B��9R��9ܐ�9�|�9�l�9FX�9H�9�;�9h1�9)�9q(�9x   x   �7�9&7�9,H�9PR�9w`�9�v�9���9
��9T��9a��9^��9���9��9���9-��9:��9[��9P��9���9��9���9u��9�u�9�`�9�Q�9�H�9I8�9�7�9V2�9m2�9x   x   I>�9�K�9(X�9r`�9o�9��9���9���9���9��9���9/��9T��9���9���9���9���94��9��9��9���9��9o�9F`�9kX�9kJ�9�=�9�>�9�:�9>�9x   x   �Y�9�a�9l�9~v�9���9e��9͞�9��9S��97��9��9|��9���9Z��9:��9���9���9y��9���9Ɵ�9���9��9�v�96l�9!b�9�Z�9�L�9�O�9tP�9M�9x   x   #m�9�p�9}�9���9���9͞�9���9|��9���9���9���9'��9,��9��9/��9���9���9��9	��9]��9���9���9�|�9�o�9�l�9ph�9�`�9�i�9`�9�h�9x   x   ��9���9ސ�9��9���9y��9x��9|��9���9��9���9���9���9���9R��9���9��93��9ح�9.��9(��9ې�9]��9��9���9x�9u�9�u�9)x�9���9x   x   2��9���9��9K��9���9S��9 ��9���92��9R��9���9���9���9���9���9��9��9���9-��9l��9��9��9��9V��9��9=��9��9<��9z��9���9x   x   ��9ҵ�9׷�9\��9��90��9���9��9V��9j��9���9
��9`��9���9`��9���9=��9M��9"��9s��9���9
��9���9��9���9���9��99��9|��9���9x   x   g��9v��9���9Y��9���9��9���9���9���9���95��9`��9v��9U��9U��99��9]��9���9��9E��9���9���9���9��9���9c��93��9K��9y��9F��9x   x   ���93��9���9���9/��9{��9&��9���9���9��9a��9���9��9���9���9���9
��9���9k��9���9��9!��9)��94��9��9���9���9W��9>��9+��9x   x   ���9b��91��9���9I��9���9+��9���9���9^��9w��9��9���9w��9���9���9@��9���9���9/��9���9I��9���9 ��9:��9���9��9���9���9y��9x   x   ���9_��9g��9���9���9Z��9��9���9���9���9Y��9���9z��9���9���9��9���9���9���9I��9v�9
�9��9�9�9O�9�
�9>�9���9/��9x   x   n��9$��9��9+��9���9<��9/��9S��9���9^��9\��9���9���9���9��9C��9���9��9��9��94�9��9��9�(�9Z �9��9�9��9��9�9x   x   ���9���9���95��9���9���9���9���9��9���9:��9���9���9��9D��9t��9��9��9��9�'�9)/�9�.�9�2�9�2�9�.�9t.�9�(�9��9L�9�9x   x   6��9��9��9_��9���9���9���9%��9��9E��9a��9��9G��9���9���9��9J�9�92�9�3�9g:�9�B�9�@�9�A�9:;�9�3�9,2�9�9s�9!�9x   x   ���95��9��9N��9<��9{��9��9;��9ù�9T��9���9���9���9���9��9��9��9�5�9RC�9�C�9FQ�9!P�9[Q�9OQ�9HC�9�B�9�6�9��9T�9��9x   x   ���9��9L��9���9��9���9��9ݭ�92��9-��9��9q��9���9���9��9��9�2�9UC�9�J�98R�9�[�9]W�9[�9�Q�9�K�9�C�9�1�9 �9��9:��9x   x   w��9Q��9C��9��9��9Ɵ�9\��93��9q��9s��9H��9���9/��9O��9��9�'�9�3�9�C�97R�9�W�97^�9�]�9�X�9R�9�B�9�3�9�(�9��9(��92��9x   x   ���9M��9S��9���9���9ƍ�9Ɛ�97��9���9���9��9��9��9~�99�9*/�9j:�9EQ�9�[�97^�9)e�9^�9�Z�9�Q�9>;�9�.�9��9��9X��9;��9x   x   ���9<��9���9u��9��9��9���9��9���9��9���92��9Q��9%
�9��9�.�9�B�9&P�9hW�9�]�9^�9�W�9�P�9�A�9�.�9O�9�	�95��9C��91��9x   x   ٛ�9���9�|�9�u�9o�9�v�9}�9g��9#��9���9���95��9���9��9��9�2�9�@�9^Q�9[�9�X�9�Z�9�P�9D@�9<3�9��9��90��9��9���9���9x   x   ̅�9q�9�l�9�`�9M`�9>l�9�o�9"��9_��9$��9��9<��9
��9�9�(�9�2�9�A�9RQ�9�Q�9R�9�Q�9�A�9=3�9�(�9�9��9��9��9r��93��9x   x   mm�9L`�9EX�9�Q�9pX�9*b�9�l�9���9��9���9���9&��9C��9��9f �9�.�9B;�9PC�9�K�9�B�9D;�9�.�9��9�9k��9���99��9v��9��9���9x   x   �Z�9-L�9H�9�H�9vJ�9�Z�9}h�9!x�9K��9ũ�9g��9���9���9Z�9��9x.�9�3�9�B�9�C�9�3�9�.�9O�9��9��9���9(��9>��9���9�x�9Fh�9x   x   $=�9�7�9�;�9O8�9�=�9�L�9�`�9#u�9��9���97��9���9��9�
�9�9�(�962�9�6�9�1�9�(�9��9�	�91��9��95��9=��9���9bu�9y`�9�L�9x   x   l7�9�2�9m1�9�7�9�>�9�O�9�i�9�u�9F��9@��9T��9g��9���9K�9��9��9�9��9# �9��9��92��9��9��9o��9}��9]u�9Fi�9�P�9Z?�9x   x   j(�9�!�9)�9[2�9�:�9�P�9`�91x�9���9���9���9H��9���9���9��9K�9s�9Y�9��9*��9\��9;��9���9q��9��9�x�9x`�9�P�979�9�2�9x   x   "�9$"�9r(�9j2�9>�9M�9�h�9���9���9���9N��95��9���9>��9#�9�9)�9��9C��9;��9>��9-��9���93��9���9@h�9�L�9X?�9�2�9�(�9x   x   k��9���9n��9x�9��9�"�9�0�9.C�9V�9[h�9+z�9���9l��9��9��9��9Ȧ�9���9���9$��9y�9/g�9�V�9B�9�1�9�$�91�9��9H��9��9x   x   ���9���9��9�
�9.�9�&�9�6�9�L�9�]�9\h�9�|�9ֈ�9G��9Ɨ�9��9=��9Օ�9���9F��9�|�9#j�9�]�9�M�956�9{%�96�9��9*�9u��9���9x   x   l��9��9��9!�9? �9�.�9�?�9"S�95^�9wq�9��9���9ȋ�9Ĕ�9���9U��9͋�9���97�9�p�9�]�95R�97@�9{0�9:�9`�9�9��9��9`��9x   x   p�9�
�9&�9�!�9�0�9�;�9�M�9�Q�9�d�9�r�9w~�9���9+��9���9���94��9���9�~�9�t�9d�9�R�9bN�9�9�9�0�9�"�9��9�
�9��9F�9��9x   x   ��9*�9? �9�0�98�9-J�9lU�9�]�9Rl�9av�9��9��9��9���9���9%��9%��9lt�9>l�9�]�9�S�9�K�9�8�9�/�9�9��9�9x�9
�9��9x   x   �"�9�&�9�.�9�;�9/J�9�O�9�\�9�i�9�t�9uy�9��9/��9��9���9V��9V�9�{�9u�9�i�9R]�9P�9�I�9�;�9�/�9�'�9#�9��9�9��9��9x   x   �0�9�6�9�?�9�M�9hU�9�\�9i�9�o�9�z�9�~�9���9���9���9G��9ć�9�}�9oy�9�p�92h�9]�9U�9�M�9?�9�6�9c0�9$+�9�&�9%�9'�95+�9x   x   .C�9�L�9$S�9�Q�9�]�9�i�9�o�9ou�9~�9*��9$��9>�9V��9Ą�9-��9�~�9#u�9�p�9�i�9?]�9TR�9�S�9M�9C�9O>�9�?�9�=�9�>�9�>�9�=�9x   x   V�9�]�9,^�9�d�9Ol�9�t�9�z�9�}�9�y�9��9��9-��9��9P~�9�y�9�~�9�y�9�t�9�l�9�d�9�\�9�]�9\V�9&T�9�L�9pN�9�Q�9�M�9PN�9=T�9x   x   Wh�9Vh�9uq�9�r�9`v�9sy�9�~�9'��9��9<��9��9���9@��9E��9���94�95z�9�u�9�r�9jr�9�i�9h�9�g�92h�9�^�9!d�9�c�9�^�9�g�9�g�9x   x   %z�9�|�9��9r~�9݀�9��9���9"��9��9��9��9ւ�9���9}��9��9��9���9b�9 �9|�9�y�9b{�9�y�9�}�9z�9�z�9E{�9�|�9kz�9~{�9x   x   }��9ˈ�9���9���9��94��9���9>�9-��9���9Ղ�9Z��9��9̓�9���9l��9=��9t��9���9���9���9���9ˍ�9H��9>��9���9��9'��9Ƌ�9���9x   x   g��9A��9���9$��9��9���9���9W��9��9D��9���9 ��9>��9c��9̋�9���9B��9Α�9���9͛�9���9���9ġ�90��9Y��9���9a��9���9q��9r��9x   x   ��9���9���9���9���9��9G��9���9U~�9N��9y��9˃�9[��9���9���9_��9o��9\��9���9ɮ�9���9q��9��9ڴ�9ϴ�9��9V��9m��9��9Z��9x   x   ���9��9���9���9���9V��9ɇ�9-��9�y�9��9��9���9ȋ�9���9���9��9���9߫�9
��9:��9��9��9���9���9r��9ѿ�9L��9
��9α�9լ�9x   x   ��9;��9T��93��9'��9X�9�}�9�~�9�~�98�9��9q��9���9d��9��90��9 ��9پ�9��9c��9���9��9��9���9)��9���9��9���9���9d��9x   x   ���9ϕ�9ϋ�9���9'��9�{�9oy�9%u�9�y�93z�9���9@��9K��9v��9���9	��9���9���9L��9i��9i��9���9���9&��9��9}��9 ��9���9���9���9x   x   ���9���9���9�~�9ot�9u�9�p�9�p�9�t�9�u�9h�9q��9Б�9[��9��9ܾ�9���90��96��9���9���9Q��9���9���9���9��9���9���9��9ު�9x   x   ���9B��95�9�t�9?l�9�i�99h�9�i�9�l�9�r�9�9��9���9���9��9��9M��98��9���91��9a��9���9���9���9���9,��9 ��9��9b��9Y��9x   x   '��9�|�9�p�9d�9�]�9Z]�9]�9D]�9�d�9lr�9|�9͈�9כ�9ˮ�9=��9g��9i��9���91��9*��9g��9���9���9���9���91��9F��9��9���9��9x   x   y�9%j�9�]�9�R�9�S�9	P�9U�9VR�9�\�9�i�9�y�9���9���9���9��9���9l��9���9f��9g��9���9K��9[��9���9���9~��9$��9\��9���9���9x   x   .g�9�]�96R�9hN�9�K�9�I�9N�9�S�9�]�9	h�9g{�9���9���9x��9
��9 ��9���9T��9���9���9J��9���9V��9���9]��9��9I��9��9ǋ�9�|�9x   x   �V�9�M�9=@�9�9�9�8�9�;�9?�9#M�9eV�9�g�9�y�9э�9̡�9��9���9 ��9���9���9���9���9Y��9S��9'��9w��9G��9ͱ�9	��9���9�y�93h�9x   x   $B�986�90�9�0�9�/�9�/�9�6�9	C�94T�9:h�9�}�9U��97��9��9���9���9*��9���9���9���9���9���9��9R��9P��9���9e��9�}�91g�98T�9x   x   �1�9�%�9?�9#�9�9�'�9j0�9S>�9 M�9�^�9z�9G��9_��9ش�9w��9/��9��9���9���9���9���9\��9K��9R��9K��9d��9�y�9�_�9�M�9%?�9x   x   �$�96�9g�9��9��9#�9.+�9�?�9rN�9$d�9�z�9���9���9���9Կ�9���9���9��91��98��9���9��9ձ�9���9e��9h|�9�c�9(N�9�>�9A)�9x   x   0�9��9!�9�
�9�9��9�&�9�=�9�Q�9�c�9W{�9���9f��9^��9N��9!��9��9���9!��9E��9��9G��9��9^��9�y�9�c�9R�9@>�9x)�9��9x   x   ��9,�9��9��9�9�9%�9�>�9�M�9�^�9�|�9-��9��9s��9��9��9���9���9��9��9^��9��9���9�}�9�_�9/N�9E>�9 #�9��9�9x   x   H��9|��9��9L�9
�9��9'�9�>�9VN�9�g�9nz�9ϋ�9z��9��9ѱ�9���9���9��9a��9���9���9ʋ�9�y�90g�9�M�9�>�9z)�9��9��9��9x   x   ���9���9c��9��9��9��9@+�9�=�9CT�9�g�9�{�9���9x��9Y��9ݬ�9n��9���9��9V��9���9���9�|�91h�90T�9#?�9C)�9��9�9��9���9x   x   ɾ�9���9��9=��9���9=��9���9��9:�9�&�9�6�9X@�9�F�9�S�9	[�9�S�9�\�9�U�9�E�9�A�9&5�9�%�9/�9��9���9��9���9;��9���9���9x   x   ���9X��9#��9Y��9���9���9 �9�	�9��9�'�9D4�9b>�9 J�9�N�9�M�9�L�9$L�9J�9P>�9I4�99)�9��9v�9k�9H��9d��9C��9 ��9���9���9x   x   !��9��9���9Z��9���9���9��9��9� �9�)�9�1�9�B�9�H�9�E�9�N�9oG�9�I�9YC�9�0�9Y)�9h �9U�9f�9h��93��9Y��9���9���9t��9X��9x   x   ?��9W��9V��9[��9���9���9b�9K�9Z&�9�/�9E1�9n@�9�@�9�E�9lD�96@�9I?�9�1�981�9�$�9a�9�9o��9Z��9���9���9���9���9��9p��9x   x   ���9���9���9���9'��9?�9[�9��9�&�9u2�9�2�9i9�9N>�9.F�9�>�9D:�9M3�9�0�9(�9��9/�9^�9���9��9���9_��92��9"��9���9L��9x   x   ;��9���9���9���9E�9��9��9��9�&�9\4�9o7�9�8�9�>�9�?�98�9�6�9�5�9d&�9��9s�9i�9�9b��9���9���9#��9��9���9���9���9x   x   ���9 �9��9\�9T�9��9�"�9x&�9�,�9G4�9t4�9?9�9A�9T8�9�5�9�2�9�,�9�&�9_"�9P�97�9��9 �9��9���9���9���9���9���9���9x   x   ��9�	�9��9J�9��9��9z&�9.�9�/�9�6�9�4�9;�9<�9�4�9{7�920�9-�9:'�9g�9r�9��9��9�	�9��9��9R�9q��9���9�9�9x   x   4�9��9� �9Z&�9�&�9�&�9�,�9�/�9�4�9�9�9�8�9~=�9�8�9d8�9�4�9�0�9s,�9�%�9�'�9�&�9��91�9Y�9F�9H�9]�9T�9{�90�9��9x   x   �&�9�'�9�)�9�/�9q2�9]4�9C4�9�6�9�9�9�5�9D:�9�8�9�7�9	;�95�9�4�9�4�9O2�9p.�9O+�9t(�9�%�9!�9�#�9� �9 �9w�9��99$�9� �9x   x   �6�9@4�9�1�9C1�9�2�9p7�9q4�9�4�9�8�9H:�9S<�9:�9�5�936�9�5�9�5�9�2�9�2�9=1�9�2�9�6�9^3�9n.�9�0�9h-�9�0�9/�910�9�.�973�9x   x   W@�9_>�9�B�9i@�9f9�9�8�979�9;�9y=�99�9:�9?�9<�9U7�99�9;�9�>�9C�9?�9�@�9�D�9�@�9�B�9<@�9�C�9 B�9�?�9C�9�@�9�D�9x   x   �F�9J�9�H�9�@�9L>�9�>�9A�9<�9�8�9�7�9�5�9<�9�@�9#@�9�<�9-A�9J�9�I�9�F�9�K�9K�9�M�9P�9cO�9�X�9)P�9zP�9	M�94K�9�L�9x   x   �S�9�N�9�E�9�E�9-F�9�?�9V8�9�4�9c8�9;�906�9]7�9'@�9F�9�E�9UE�9�M�9T�9LS�9\�9"]�9,a�9e�9�`�92a�9d�9a�9^�9�Z�9�R�9x   x   [�9�M�9�N�9jD�9�>�98�9�5�9y7�9�4�95�9�5�99�9�<�9�E�9�N�9�M�9C\�9_�91a�9l�9�k�9�q�9+u�9�j�9�t�9"s�9Ok�9�k�9}b�9`�9x   x   �S�9�L�9qG�95@�9F:�9�6�9�2�910�9�0�9�4�9�5�9;�9)A�9SE�9�M�9S�9�[�9�f�9�n�9�p�9t�9�{�9~�90~�9�{�9�s�9Cq�9�n�9�d�9E\�9x   x   �\�9%L�9�I�9A?�9P3�9�5�9�,�9-�9x,�9�4�9�2�9�>�9�I�9�M�9B\�9�[�9sd�9t�9�{�9w��9h��9|��9|��9σ�9L��9���92{�9du�9e�9[�9x   x   �U�9J�9_C�9�1�9�0�9k&�9�&�9='�9�%�9Q2�9�2�9
C�9�I�9"T�9_�9�f�9t�9 |�9F��9M��9E��9ې�94��9A��9���9C��9{�9�s�9�f�9�]�9x   x   �E�9M>�9�0�961�9(�9��9["�9h�9�'�9p.�9D1�9?�9�F�9RS�94a�9�n�9�{�9F��9���9M��9��9��9���9���9\��9���9�{�91n�9c�9)R�9x   x   �A�9E4�9Z)�9�$�9��9w�9V�9u�9�&�9S+�9�2�9�@�9�K�9\�9	l�9�p�9|��9N��9I��9���9̗�9���9v��9��9��9ɀ�9*r�9hj�97\�9KL�9x   x   %5�9<)�9i �9d�9/�9j�9?�9��9��9}(�9�6�9�D�9K�9(]�9�k�9#t�9k��9I��9 ��9˗�9|��9ɗ�9���9��9��9�r�9�l�9L]�9�J�9OD�9x   x   �%�9��9U�9�9g�9�9��9��92�9�%�9j3�9�@�9�M�92a�9�q�9�{�9y��9ڐ�9��9���9ŗ�9ș�9;��9���9�|�9r�9�a�9�M�9�@�9�4�9x   x   )�9w�9b�9q��9���9c��9 �9�	�9]�9!�9{.�9�B�9P�9e�93u�9~�9���9:��9���9y��9���9@��9���9�}�9�u�9�c�9�O�9	C�9 -�9p!�9x   x   ��9k�9j��9^��9��9���9��9��9O�9�#�9�0�9<@�9iO�9�`�9�j�93~�9҃�9K��9���9��9��9���9�}�96j�9,a�9�P�9�?�92�9�#�9E�9x   x   ���9N��96��9���9���9���9���9��9S�9� �9j-�9�C�9�X�92a�9�t�9�{�9H��9}��9\��9���9��9�|�9�u�9$a�9wW�9�B�9�,�9� �9�9�9x   x   ��9e��9V��9���9`��9(��9��9Y�9h�9
 �9�0�9B�91P�9d�9(s�9�s�9ǁ�9J��9���9ɀ�9�r�9!r�9�c�9�P�9�B�9�2�9 �9+�97�9���9x   x   ���9F��9���9���95��9$��9���9v��9Z�9z�9/�9�?�9�P�9a�9Tk�9Eq�95{�9{�9�{�9-r�9�l�9�a�9�O�9�?�9�,�9�9��9Q��9���9b��9x   x   A��9��9���9���9%��9���9��9���9�9 �9;0�9C�9M�9^�9�k�9�n�9ju�9�s�94n�9oj�9M]�9�M�9C�92�9� �9$�9N��9���9���9i��9x   x   ���9���9v��9��9���9���9���9�99�9=$�9�.�9�@�98K�9�Z�9�b�9�d�9 e�9�f�9c�9?\�9�J�9�@�9-�9�#�9�93�9���9���9���9���9x   x   ���9���9U��9v��9T��9���9���9�9��9� �9<3�9�D�9�L�9�R�9`�9C\�9[�9�]�9.R�9OL�9ND�9�4�9m!�9K�9�9���9c��9k��9���9���9x   x   ��9���9��9`��9��9ʱ�9ݻ�9!��9���9���9R��9*��9� �9��9��9�9��9��9I �9���9���9���9���9���9���9��9��9@��9��9&��9x   x   ڒ�9���9���9���9ũ�9��9۸�9���9~��9!��9f��9��9���9��9��9��9� �9���9���9���9��98��9���97��9h��9#��9��9���9���9��9x   x   ��9���9��9��9Z��9���9���9���9���9���9b��9P��9H��9 �9���9p �9V��9���9��9��9]��9���97��9��9���9��9v��9���9���9��9x   x   c��9���9��9z��9��9r��9<��9���9T��9��9��9��9X��9-��9a��9{��9���9���9���9��9���9���9���9���9��9���9��9���9>��9˝�9x   x   ��9ĩ�9^��9
��9���9k��9J��9T��9��9Z��9���9N��9���9���9O��9y��9��9i��9O��9��9���9���9~��9���9���9���9_��9T��9��91��9x   x   Ǳ�9��9���9k��9l��9���9���9���9 ��9���9���9���9���9��9N��9���9���9��9���92��90��9���9e��9H��9R��9`��9��9r��9���9w��9x   x   ڻ�9ݸ�9���99��9O��9���9���93��9���9���9��9���9y��9D��9���9���9���9��9S��9���9��9��9)��9V��9ٻ�9��9)��9���9X��9ָ�9x   x   ��9���9���9���9Q��9���90��9R��9h��9M��9���9���9��9���9���9���93��9d��9���9���9b��9B��9���9���9[��9���9���9��9���9���9x   x   ���9z��9���9Q��9��9��9���9r��9���9D��9���9��9���9a��9���9���9���9|��9���9���9���9J��9���9P��9���9���9c��9���9���9h��9x   x   ���9"��9���9��9X��9���9���9M��9D��9���9��9N��9���9��9R��9���9^��9i��9���9���9���9���9���9��9-��9���9���9P��9 ��9���9x   x   I��9b��9b��9��9���9���9��9���9���9��9���9���9���9���9x��9N��9g��9 ��9���9���9���9���9���9���9%��9��9��9���9��9���9x   x   &��9��9J��9��9L��9���9���9���9��9M��9���9&��91��9���9���9���9���9���90��9~��9R��9{��9���9���9"��9���9���9���9���9;��9x   x   � �9���9>��9T��9���9���9y��9��9���9���9���9-��9j��9(��9���9���9���9A��9� �9� �9��9�9��9�9��9��9�9��9$�9��9x   x   ��9��9 �9,��9���9��9B��9���9a��9��9���9���9%��93��9���9���9��9��9�	�9�9��9+�9��9��9��9��9�9��9{�9?	�9x   x   ��9��9���9`��9K��9P��9���9���9���9U��9y��9���9���9���9���94�9I�9��9l�9�9;�9o�9�9�!�9�9��9z�9��9��9T�9x   x   �9��9l �9z��9y��9���9���9���9���9���9N��9���9���9���9>�9&�9M�9\�9��90!�9G(�9I&�9o(�98(�9U%�9�(�9� �9e�9��9��9x   x   ��9� �9S��9���9��9���9���97��9���9c��9i��9���9���9��9K�9M�9_�9N�9#�9�(�9�/�9�0�9�,�9�1�91/�9y)�9�#�9c�9��9/�9x   x   ��9{��9���9���9k��9��9��9j��9x��9l��9���9���9G��9��9��9Z�9T�9�#�9�-�991�9>�9�9�98�9n>�9�0�9q-�9�"�9��9�9g�9x   x   K �9���9��9���9V��9���9V��9���9���9���9���94��9� �9�	�9q�9��9#�9�-�940�9�7�9�<�9�7�9R=�9�7�9�0�9�.�9�#�9��9�9<	�9x   x   ���9���9��9��9��96��9���9���9���9���9���9���9� �9�9�95!�9�(�9<1�9�7�9W:�9�?�9h@�9s9�98�90�9(�93"�9�9��9� �9x   x   ���9��9^��9���9���92��9��9f��9���9���9���9W��9��9��9>�9F(�9�/�9>�9�<�9�?�9�N�9	@�9v=�9d>�9�1�9�&�9n�9��9��9l��9x   x   ���98��9���9���9���9���9��9G��9O��9���9���9~��9�9.�9q�9M&�9�0�9�9�98�9p@�9@�9�7�9�8�9-/�9�&�9G�9��9��9��9s��9x   x   ���9���9>��9���9���9j��9.��9���9���9���9���9���9��9��9�9u(�9�,�98�9K=�9u9�9t=�9�8�93/�9�'�9��9�9?�9C��9H��9���9x   x   ���9=��9��9���9���9N��9Y��9���9S��9��9���9���9�9��9�!�95(�9�1�9q>�9�7�98�9d>�9(/�9�'�9�"�9��9�95��9m��9���9R��9x   x   ���9a��9���9��9���9P��9ۻ�9]��9���93��9*��9/��9��9��9#�9\%�98/�9�0�9�0�90�9�1�9�&�9��9��9B�9���9.��9(��9���9>��9x   x   ��9&��9��9���9��9c��9��9��9���9���9��9���9��9��9��9�(�9~)�9p-�9�.�9(�9�&�9I�9�9�9���9/��9���9���9̺�9w��9x   x   ��9��9y��9��9b��9��9,��9���9f��9���9��9���9�9�9}�9� �9�#�9�"�9�#�93"�9n�9��9>�98��9*��9���9��9���9@��9���9x   x   D��9���9�9���9V��9x��9���9��9���9W��9���9���9��9��9��9e�9d�9��9��9�9��9��9A��9m��9+��9���9���9��9��9H��9x   x   ��9���9���9C��9	��9���9]��9���9���9��9��9���9(�9y�9��9��9��9�9�9��9��9��9L��9���9���9Ѻ�9A��9��9ʢ�9���9x   x   (��9��9��9Ν�97��9���9ظ�9���9d��9���9���9A��9��9A	�9Y�9��94�9m�9=	�9� �9n��9s��9���9N��9=��9w��9���9I��9���9]��9x   x   �U�9v]�9:a�9e�9�p�9�w�9�{�9L��9$��9r��9���9h��9'��9x��99��9���90��9H��9���9���9H��9P��9Ő�9���9|�9�w�94q�9,d�9�c�9�]�9x   x   v]�9P_�93c�9d�9�m�9�z�9V��9���9��9��9/��9��9c��9���9���9��9���9ϵ�9���9���9��9��9a��9���9�y�9El�9ie�9�a�9�]�9�^�9x   x   9a�98c�9=l�9�i�9Tv�9|�9���9l��9���9���9է�9f��9���9J��9)��9b��9S��9+��9���9���9ژ�9���9��9|�9Ox�9Pi�9�l�9�d�9�`�9�`�9x   x   e�9d�9�i�9�u�9�z�9��9u��9��9���9��9���95��9+��9���9x��9	��9B��9��9ۢ�9כ�9ӓ�9���9���9�x�9�u�9%i�9[c�9xe�9{_�9`�9x   x   �p�9�m�9Pv�9�z�9�~�9���9���9t��9���9}��9֦�9���9*��9ܯ�9!��9��9���9���9ĝ�9��9���9A��9��9�z�9w�9-o�9�o�9�m�94i�9�l�9x   x   �w�9�z�9|�9��9���9��9v��9r��9��9���9���9��9��9��9ƪ�9��9p��9��9���9���9Ҕ�9?��9��9|�9�x�9�w�9nt�9�p�9�q�94t�9x   x   �{�9N��9���9q��9}��9w��9��9H��9���9���9ѧ�9k��9���9���9��9w��9���9Ϛ�9L��9���9P��9b��9���9���9 |�9�z�9z�9�x�9z�9=z�9x   x   I��9��9i��9��9n��9p��9E��9-��9r��98��9b��9Ĩ�9b��9
��9=��9x��9t��9��9ߝ�9T��9-��9���9}��9��9E��9=��9e��9���9���9"��9x   x   $��9ݒ�9���9���9���9��9���9p��9Ƣ�9)��9!��9Z��9���9&��9���9���9���9��9��9��9"��9��9���9��9���9��9��9#��9���99��9x   x   m��9��9���9|��9z��9���9���96��9+��9��9��9���9��9A��9��9q��9���9 �9���9&��9��9��9��9��9J��9/��9c��9���9���9���9x   x   ���9+��9Ч�9���9Ԧ�9���9ҧ�9^��9!��9��9h��9��95��9y��9
��9y��9T��9���9���9���9���9Ħ�9��9��9���9��9-��9s��9Z��9���9x   x   e��9���9e��9<��9}��9��9j��9ɨ�9]��9���9��9k��9���9���9��9ϭ�9��9���9~��9���9F��9ɪ�9>��9��9
��9+��9���9��9���9��9x   x   #��9c��9���9+��9'��9��9���9e��9­�9��97��9���9S��9���9��9Ҳ�9��9���9}��9��9��9۶�9J��94��9ɶ�9Ѻ�9���93��9���9���9x   x   u��9���9D��9���9د�9��9���9��9(��9C��9z��9���9���9X��9��9���9���9���9��9l��9D��9���9���9g��9���9T��9���9���9��9��9x   x   7��9���9+��9z��9��9ɪ�9��99��9���9��9��9��9���9��9`��9���9��9K��9p��9e��9���9���9���9��9���9��9���9���9���9��9x   x   ���9��9[��9��9��9��9w��9x��9���9t��9y��9Э�9ղ�9���9���9���9���9��9$��9a��9���98��9"��91��9���9L��9���9Q��9���98��9x   x   .��9���9X��9F��9���9v��9���9s��9���9���9X��9��9!��9���9��9���9#��9S��9b��9e��9���9���9���9C��9c��9��9���9���9��9���9x   x   D��9ε�9)��9��9���9��9К�9��9��9Ġ�9���9���9���9���9O��9��9V��9���9��9���9e��9���9q��9���9���9I��9���9=��9��9���9x   x   ���9���9���9ޢ�9ŝ�9���9P��9��9	��9���9���9~��9~��9��9s��9��9c��9��9��9���9���9s��9���9���9D��9C��9���9��9���99��9x   x   ���9���9���9֛�9��9���9���9V��9��9)��9��9���9��9n��9g��9e��9g��9���9���9]��9��9���9���9��9���9��9O��9���9^��9���9x   x   E��9��9ߘ�9ӓ�9���9Ք�9T��90��9'��9��9���9G��9���9C��9���9���9���9k��9���9��9@��9G��9���9<��9���9���9���9���9���9���9x   x   Q��9��9���9���9D��9D��9d��9Ð�9��9��9Ȧ�9ͪ�9��9���9���9=��9���9���9z��9���9E��9q��91��9i��9��9
��9���9ȷ�9l��9��9x   x   Ȑ�9Y��9��9���9��9��9���9z��9���9��9!��9>��9K��9���9���9$��9���9q��9���9���9���95��9���9K��9)��9K��9��9w��9���9ɚ�9x   x   ���9���9|�9�x�9�z�9|�9��9��9��9���9��9	��96��9p��9��9,��9I��9���9���9��9:��9l��9I��9���9���9���9߯�9���9כ�9���9x   x   |�9�y�9Px�9�u�9w�9�x�9	|�9F��9���9M��9���9��9ȶ�9���9���9���9g��9���9L��9���9���9��9'��9���9��9���9$��9���9���9��9x   x   �w�9Il�9Ti�9)i�97o�9�w�9�z�9G��9��93��9��9-��9պ�9T��9��9O��9��9E��9A��9��9���9��9H��9���9���9Ȥ�9J��9Ώ�9"��9�y�9x   x   2q�9ie�9�l�9Wc�9�o�9kt�9z�9k��9��9l��94��9���9���9���9���9���9���9���9���9P��9���9���9��9��9(��9M��9v��9o��9Lz�9ht�9x   x   .d�9�a�9�d�9ze�9�m�9�p�9�x�9���9 ��9���9w��9��98��9���9���9S��9���9?��9��9���9���9̷�9t��9���9���9̏�9m��9�y�9q�9�l�9x   x   �c�9�]�9�`�9}_�97i�9�q�9z�9��9���9���9^��9��9���9!��9���9���9 ��9��9���9`��9���9l��9���9ԛ�9���9��9Lz�9�p�9*j�9�_�9x   x   �]�9�^�9�`�9
`�9�l�90t�9@z�9&��9A��9ǚ�9���9~��9 ��9��9��9;��9���9���95��9���9���9��9̚�9���9��9�y�9ft�9�l�9�_�9�^�9x   x   �!�9_&�9&*�9u+�9�2�9y4�9B�9QH�9�P�9hZ�9d�9bh�9�h�93s�9�y�9�s�9�x�9jr�9i�9[i�9�d�92[�9�O�9�G�9�A�9�3�9S3�9�*�9�,�9�&�9x   x   `&�9,�9�'�9�2�9�6�9
>�9�H�9�I�9DU�9GZ�92`�9yh�9�m�9�o�9p�9Iq�9�o�9jn�9�g�9�^�9gY�9V�9�J�9VH�9�>�9�5�9�3�9�&�9G*�9�&�9x   x   %*�9�'�9�1�9�5�9�7�9�?�9�B�9�K�9�U�9�Y�9�]�9ej�9�k�9�i�9Bo�9�h�9�k�9j�9&_�9�[�9%U�9�J�9C�9�?�9/8�9V5�9?2�9�(�9 +�9Z)�9x   x   q+�9�2�9�5�9Z6�9A�9�E�9HM�9�R�9T[�91_�9J^�9�h�9wg�9Bl�9�l�9dh�9mh�93^�9D]�9�Z�9�S�9zM�9 F�9�?�987�95�9G2�9'+�9�,�9.�9x   x   �2�9�6�9�7�9A�9�E�97I�9:R�9�S�9LZ�9�a�9d�9�f�9e�9�d�9�d�9f�9�d�9�b�9w[�9JS�9�Q�9$H�9(G�9�@�9D7�9R8�9�2�9:.�9D1�9�-�9x   x   y4�9>�9�?�9�E�99I�9�J�9�T�9�W�9�\�9�d�9�d�9�e�9Ti�9>i�9�e�9�d�9]c�9�\�9LW�9qT�9�L�9IH�9 E�90@�9,=�9�3�9o3�9�6�9�6�93�9x   x   B�9�H�9�B�9FM�96R�9�T�9;]�95`�9�^�9Cb�9�c�9�c�9hj�9Gd�9�c�9�b�9�_�9�_�9�^�9�R�9oR�9�M�9�B�9�I�9ZB�9�<�9@�9�8�9<A�9<<�9x   x   SH�9�I�9�K�9�R�9�S�9 X�97`�9�b�9�_�9�e�9�c�9Eg�9tf�9.c�9�e�9_�9�b�9�_�9JX�9�S�9R�9�K�9�H�9�G�9UE�9�E�96@�9�>�9
F�9WE�9x   x   �P�9CU�9�U�9V[�9GZ�9�\�9�^�9�_�9?g�9.h�9�b�9<e�9�c�9�h�9�g�9�_�9�_�94[�99[�9�[�9$U�9>V�9�Q�9�Q�9�N�9�J�9O�9�J�9+O�9�Q�9x   x   fZ�9EZ�9�Y�94_�9�a�9�d�9Db�9�e�92h�9�b�9-d�9 d�9�a�9wg�9�f�9>a�9�e�9ob�9 ]�9+[�9|Y�9^Y�9�V�9DY�9aX�9%Z�9g[�9�W�9Y�9�V�9x   x   d�92`�9�]�9H^�9d�9�d�9�c�9�c�9�b�91d�9�l�9Od�9�d�9:c�9Ud�9d�9ac�9�_�9j^�9�_�9we�9I`�9�\�9_�9�_�9�_�9�^�9�_�9�\�92`�9x   x   _h�9{h�9]j�9�h�9�f�9�e�9�c�9Dg�96e�9&d�9Ud�99d�9�f�9-c�9af�9jg�9�g�9j�9�g�9*h�9�k�9�g�9�m�9�f�9�j�9Rj�9�g�9am�9�g�9dl�9x   x   �h�9�m�9�k�9vg�9e�9Zi�9jj�9vf�9�c�9�a�9�d�9�f�9l�9�h�9kc�9�h�9�k�9|n�9<j�9o�9o�9�r�9:s�9|p�9-v�9�p�9Vr�9t�9!n�9�o�9x   x   -s�9�o�9�i�9<l�9�d�9Bi�9Id�9/c�9�h�9tg�9:c�92c�9�h�9Fg�9�k�9�h�9To�9�q�9q�9�v�9�x�9y�9�}�9h{�9U{�9�}�9�x�9�x�9Nv�9lq�9x   x   �y�9p�9?o�9�l�9�d�9�e�9�c�9�e�9�g�9�f�9Vd�9`f�9kc�9�k�9�o�9�p�9�z�9}�9�{�9���9�~�9���9��9=}�9׃�91��9�}�9���9U{�9V|�9x   x   �s�9Gq�9�h�9bh�9f�9�d�9�b�9_�9�_�9=a�9d�9jg�9�h�9�h�9�p�9Rr�9�w�9g|�9*��9��9I��9��9އ�9���9���9<��95��9ˀ�9�}�9x�9x   x   �x�9�o�9�k�9ch�9�d�9]c�9�_�9�b�9�_�9�e�9dc�9�g�9�k�9[o�9�z�9�w�9�z�9��9e��9S��9���9y��9(��9ԏ�9\��9���9���9Y��9�y�9�w�9x   x   gr�9nn�9j�99^�9�b�9�\�9�_�9�_�9=[�9nb�9�_�9j�9�n�9�q�9}�9f|�9��9��9G��9O��9���9���91��9?��9���9���9J��9��9<}�9�}�9x   x   i�9�g�9+_�9E]�9u[�9OW�9�^�9HX�9=[�9]�9o^�9�g�9>j�9q�9�{�9.��9g��9H��9��9\��9ѓ�9��9ޕ�9���9	��9���9V��9��9}z�9bq�9x   x   Xi�9�^�9�[�9�Z�9NS�9tT�9�R�9�S�9�[�9+[�9�_�9(h�9o�9�v�9���9��9U��9L��9V��9��9Z��92��9��9˒�9'��9��9���9���9w�9�n�9x   x   �d�9fY�9&U�9�S�9�Q�9�L�9pR�9R�9(U�9Y�9|e�9�k�9o�9�x�9�~�9J��9���9���9ד�9Z��9���9���9V��9��9
��9��9�}�9ux�9�n�9�k�9x   x   2[�9V�9�J�9�M�9)H�9MH�9�M�9�K�9BV�9_Y�9T`�9�g�9�r�9y�9���9$��9w��9���9��93��9���9���9��9_��9���9���9�y�9�s�93h�9O_�9x   x   �O�9�J�9C�9"F�9&G�9E�9�B�9�H�9�Q�9�V�9�\�9�m�9=s�9�}�9��9��9.��93��9��9��9Y��9��9��9u��9��9}�9mr�9Xm�9Q]�9eV�9x   x   �G�9ZH�9�?�9�?�9�@�90@�9�I�9�G�9�Q�9AY�9_�9�f�9}p�9p{�9A}�9���9Տ�9?��9���9˒�9��9a��9x��99~�9�z�9Yq�9ng�9�^�9�Y�9lR�9x   x   �A�9�>�9.8�9<7�9J7�9/=�9`B�9QE�9�N�9iX�9�_�9�j�93v�9V{�9ڃ�9���9Y��9���9��9(��9��9���9��9�z�9nv�9�i�9�_�9oW�9�M�9F�9x   x   �3�9�5�9S5�95�9S8�9�3�9�<�9�E�9�J�9-Z�9�_�9[j�9�p�9�}�93��9D��9��9���9�9��9��9Ą�9}�9Zq�9�i�9�_�9�Z�9�L�9E�9�<�9x   x   S3�9�3�9D2�9I2�9�2�9n3�9@�98@�9O�9j[�9�^�9�g�9\r�9�x�9�}�98��9���9N��9T��9���9�}�9�y�9lr�9qg�9�_�9�Z�99M�9�?�9�@�9�3�9x   x   �*�9�&�9�(�9(+�9<.�9�6�9�8�9�>�9�J�9�W�9�_�9hm�9t�9�x�9���9̀�9Z��9��9��9���9nx�9�s�9Wm�9�^�9pW�9�L�9�?�9Q9�9�5�9;-�9x   x   �,�9C*�9#+�9�,�9D1�9�6�9BA�9F�91O�9Y�9�\�9�g�9n�9Vv�9X{�9�}�9�y�9>}�9�z�9w�9�n�95h�9R]�9�Y�9�M�9E�9�@�9�5�93�9-�9x   x   �&�9�&�9^)�9.�9�-�93�9C<�9WE�9�Q�9�V�95`�9cl�9�o�9oq�9O|�9x�9�w�9�}�9bq�9�n�9�k�9J_�9eV�9pR�9F�9�<�9�3�9<-�9-�9�'�9x   x   ���9���9���90��9���9� �9��9��9��9��9��9�"�9�+�9M)�9�,�9z-�9�+�9�(�9�,�9�"�9��9k�9��9&	�9��9���9[��9 ��9���9���9x   x   ���9)��9��9r��9���9���9��96�9�91�9�#�9&�9�#�9_)�9�-�9E.�9*�9�#�9X%�9u#�9�9��9+
�9��9���9���9��9��9��9}��9x   x   ���9
��9+��9���9���9��9Z
�9v�9�9��9�#�9� �9}&�9j(�9�(�9�'�9N&�9� �9�$�9��9��9��9��9{�9���9f��9'��9v��9���9���9x   x   2��9n��9���9���9���9��9(�9��9��9��9��9�"�96&�9(�9I(�9�&�9�"�9|�9��9k�9O�9m�9��9J��9���9J��9]��9���9���9���9x   x   ���9���9���9���9��9�9X�9��9#�9��9��9A#�9�&�9%�9�&�9�"�9��9~�9��9��9k�9Z�9��92��9���9���9���9���9b��9���9x   x   � �9���9��9��9�9_�9{�9��9��9h�9� �9p%�9C �9��9�%�9
!�9��9��9��9p�9��9�9[�9%�9���9~��9W��9���9���9���9x   x   ��9��9Y
�9&�9X�9y�9��9��9�9K�9%�9� �9��90!�9b$�9��9)�9��9�9�9X�9�9�
�9��9(�9��96�9��9��9��9x   x   ��93�9w�9��9��9��9��9��9��9��9�!�9I#�9�"�9�!�9��9��9�9��9��9��9��9��9"
�9��9��9��9�
�9�9�9��9x   x   ��9�9�9��9#�9��9�9��9��9��9� �9��9!�9��9N�9�9S�9+�9Q�9��9��9��9��9��9I�9?�9Z�91�9��9�9x   x   ��93�9��9��9��9b�9J�9��9��9l#�9!�9�!�9f"�9\�9��9�9Y�9/�9%�9�9��9��92�9��9��9f�9��92�9{�9��9x   x   ��9�#�9�#�9��9��9} �9%�9�!�9� �9!�9
$�9*!�98"�9
!�9V%�9� �9��9��9 $�9�#�9��9��9g�9��9��9M�9��93�9��9��9x   x   �"�9&�9� �9�"�9D#�9r%�9� �9J#�9��9�!�9)!�9�9�"�9r �9�%�9
#�9�"�9*!�9G%�9�!�9� �9(�9i&�9�&�9�$�9$�9�&�9q&�9J'�96!�9x   x   �+�9�#�9~&�96&�9�&�9A �9��9�"�9!�9d"�99"�9�"�9��9��9�&�9�&�9�%�9�#�9-�9�.�9y(�9�+�9�+�9�+�9 -�9�,�9+�9a,�9�(�9v.�9x   x   M)�9\)�9l(�9(�9%�9��9+!�9�!�9��9b�9	!�9m �9��9&�9�'�9�(�9�)�9#(�9�/�9�/�9/�9�/�9H/�9�3�9@3�9�.�9�/�9/�9q/�9�0�9x   x   �,�9�-�9�(�9I(�9�&�9�%�9e$�9��9M�9��9X%�9�%�9�&�9�'�9)�9�-�9-�9�-�9�/�9C5�9�:�9R8�9�8�9o?�9�8�9m9�9:�9(5�9�/�9�,�9x   x   {-�9G.�9�'�9�&�9�"�9!�9��9��9|�9!�9� �9#�9�&�9�(�9�-�9-�9�3�9v9�9V9�9;�9w@�9.?�9$B�9�B�9C>�9�?�9�;�9�9�9�9�9�3�9x   x   �+�9*�9N&�9�"�9��9��9%�9�9P�9U�9��9�"�9�%�9�)�9-�9�3�9�:�9*;�9�<�9z@�9�C�9E�9�@�9�E�9]D�9�@�9�;�9D:�9Y;�9�4�9x   x   �(�9�#�9� �9|�9�9��9��9��9.�90�9��9*!�9�#�9 (�9�-�9w9�9);�9�=�9C�9�C�9�L�9I�9�G�9 L�9�C�9C�9g?�9c;�9>8�9.�9x   x   �,�9R%�9�$�9��9��9��9�9��9S�9(�9�#�9J%�9-�9�/�9�/�9W9�9�<�9C�9�@�9kI�9�G�9�D�9<I�9dI�9,A�9 B�9�;�9\:�9�/�9�/�9x   x   �"�9y#�9��9o�9��9s�9�9��9��9�9�#�9�!�9�.�9�/�9E5�9;�9z@�9�C�9dI�9�H�9�J�9J�9	H�9GI�9|D�9�A�9�:�9Y5�9�/�9U.�9x   x   ��9�9��9M�9o�9��9X�9��9��9��9��9� �9|(�9/�9�:�9y@�9�C�9�L�9�G�9�J�9sX�9�J�9�H�9L�9�B�9A�9::�9�.�9!)�9� �9x   x   h�9��9��9k�9[�9	�9�9��9��9��9��9(�9�+�9�/�9V8�91?�9E�9I�9�D�9J�9�J�9RD�9H�9�F�9j>�9N8�9t0�9�+�9�'�9��9x   x   ��91
�9��9��9��9b�9�
�9*
�9��92�9n�9l&�9�+�9M/�9�8�9#B�9�@�9�G�96I�9	H�9�H�9xH�9�?�9BB�9�9�9�.�97+�9X&�9��9��9x   x   '	�9��9z�9O��94��9%�9��9��9��9��9��9�&�9�+�9�3�9n?�9�B�9�E�9	L�9eI�9NI�9L�9�F�9BB�9�>�9v3�9O,�9'�9��9��9��9x   x   ��9���9���9���9���9���9*�9��9O�9��9��9�$�9 -�9?3�9�8�9G>�9`D�9�C�9(A�9�D�9�B�9k>�9�9�9x3�9%-�9$�92�9��9��9>�9x   x   ���9���9k��9M��9���9���9��9��9>�9e�9R�9$�9�,�9�.�9l9�9�?�9�@�9!C�9B�9�A�9�@�9J8�9�.�9Q,�9$�9��9y�9�9s�9��9x   x   ^��9��9-��9`��9���9^��9<�9�
�9Z�9��9��9�&�9+�9�/�9:�9�;�9�;�9f?�9�;�9�:�98:�9t0�93+�9'�91�9v�9��9�
�9��9���9x   x   #��9y��9v��9���9���9���9��9#�96�97�9<�9u&�9a,�9)/�9*5�9�9�9D:�9f;�9]:�9Z5�9�.�9�+�9X&�9��9��9�9�
�9��9���9���9x   x   ��9��9���9���9c��9���9��9�9��9z�9��9M'�9�(�9s/�9�/�9�9�9Z;�9B8�9�/�9�/�9!)�9�'�9��9��9��9t�9��9���9���9���9x   x   ���9z��9���9���9���9���9��9��9��9��9��9:!�9v.�9�0�9�,�9�3�9�4�9.�9�/�9R.�9� �9��9��9��99�9��9���9���9���9���9x   x   ���9��9
��9ط�9g��9���9��9���9x��9���9k��9[��9���9r��9>��97��9���9���9p��9���9���9-��9���9��9��9���94��9"��9Y��9���9x   x    ��9;��9��9���9��9W��9���9��9���9��9��9���9q��9���9��9m��9���9r��9���97��9���9���9m��9���9���9Ҿ�9j��9��9���9��9x   x   ��9��9[��9��9���9���9���9~��9���9���9
��9���9t��9���99��9U��9��9l��9���9P��9��9���9~��9���9=��9ҽ�9���9���9���9ȼ�9x   x   ݷ�9���9��9��9���9y��9f��9��9���9���9<��9���9X��9���9���9I��9d��9r��9���9��9?��9���9I��9%��9/��9½�9߸�9��9���9��9x   x   d��9��9���9���9}��9k��9���9���9���9���9���9���9q��9D��9���9+��9���9z��9���9���9���9���9-��9!��9��9��9d��9���9x��9��9x   x   ���9U��9���9y��9l��9���9���9;��9{��9���9���9;��9���9��9h��9-��9S��9���9��9���9t��9��9���9��9���9���9��9u��9V��9 ��9x   x   ��9���9���9f��9���9���9���9��9���9��9E��9���9&��9@��9��9H��9���9��9���9���94��9���9?��9���9��9���9���9���9ټ�9a��9x   x   ���9��9{��9 ��9���9;��9��9���9j��9 ��9B��9r��9^��9v��9���9���9,��9���9%��9Z��90��9��9h��9���9���9���9>��9���9F��9��9x   x   }��9���9���9���9���9���9���9i��9���9���9���9r��9g��9A��9C��9���9h��9N��9���9W��9���9g��9���9���9f��9��9	��9���9���9���9x   x   ���9��9���9���9���9���9��9��9���9���9���9h��9O��9K��9?��9���9o��9���9<��9���9���9���9���9���9`��9X��9Z��9���9���9���9x   x   m��9��9��98��9���9���9E��9C��9���9���9y��9���9���9q��9k��9��9���9���9���9���9:��9���9r��9n��9��9���9���9���9��9N��9x   x   [��9���9���9���9���9:��9���9v��9t��9c��9���9���9z��9���9���9���96��9z��9���9���9���9[��9��9���9���9���9���9���9Z��9T��9x   x   ���9l��9t��9U��9l��9���9$��9a��9m��9O��9���9z��9e��9\��9,��9#��9M��9���9<��9���9���9c��9���9c��9��9 ��9��9���9���9���9x   x   u��9���9���9���9J��9��9C��9t��9A��9J��9n��9��9e��9:��9J��9���9���9p��9#��9���9E��92��9���9���9��9���9���9���9s��9���9x   x   B��9��95��9���9���9j��9��9���9>��9;��9i��9���9.��9E��9v��9���9p��9���9���9���9
��9W��97��9��9=��9j��9a��9���9K��9m��9x   x   5��9h��9P��9E��9&��9+��9I��9���9���9���9��9���9"��9���9���9���9���92��9C��9��9$��9���9���9���9h��9��9d��9��9`��9���9x   x   ���9���9	��9d��9���9X��9���90��9j��9r��9���97��9P��9���9o��9���9���9x��9���9���9���9(��9���9P��9:��9��9r��9���9g��9���9x   x   ���9s��9t��9n��9}��9���9��9���9O��9���9���9~��9���9s��9���91��9y��9���9���90��9���9��9���9*��9���9"��9D��9K��9p��9���9x   x   q��9���9���9���9���9��9���9#��9���9A��9���9 ��9@��9(��9���9B��9���9���9�9
�9u�96�9-�9� �9v�9���9���9���9��9���9x   x   ���95��9S��9��9���9���9���9Z��9Q��9���9���9���9���9���9���9
��9���93��9�9?��95�9� �9 �9\�9��9a��94��9���9��9���9x   x   ���9���9��9D��9���9r��99��9:��9���9���97��9���9���9D��9
��9&��9���9���9s�98�9� �95�9��9��9���9}��9*��9���9p��9���9x   x   /��9���9���9���9���9��9���9��9j��9���9���9_��9h��9/��9X��9���9&��9��97�9� �97�9J�9��9���9���9��9z��9���9z��9
��9x   x   ���9j��9���9I��9-��9���9@��9f��9���9���9u��9��9���9���9;��9���9���9���9/�9 �9��9��9��9.��9���9j��9j��9N��9���9���9x   x   ��9���9���9%��9 ��9��9���9���9���9���9r��9���9h��9���9	��9���9Q��9'��9� �9\�9��9���9+��9L��9���9a��9{��9���9���9���9x   x   ��9���9:��9-��9��9���9��9���9h��9b��9���9���9��9��9=��9m��9<��9���9w�9��9���9���9���9���9c��9���9���9���9���9W��9x   x   ���9־�9Խ�9���9��9���9���9���9��9]��9���9���9��9���9k��9��9��9%��9���9^��9}��9��9h��9a��9���9��9���9���9���9���9x   x   2��9j��9���9߸�9e��9��9���9B��9��9b��9���9���9��9���9g��9h��9u��9G��9���93��9/��9z��9l��9~��9���9���9���9���9���9���9x   x   $��9��9���9��9���9u��9���9���9���9���9���9���9 ��9���9���9#��9���9K��9���9���9���9���9O��9���9���9���9���9M��9���9߽�9x   x   Z��9��9���9���9{��9V��9޼�9L��9���9���9��9W��9���9r��9K��9\��9b��9q��9��9��9l��9r��9���9���9���9���9���9���9��9���9x   x   ��9��9ż�9��9��9 ��9c��9��9���9���9M��9V��9���9���9u��9���9���9���9���9���9���9��9���9���9X��9���9���9��9���9��9x   x   s�9,}�9�{�9��9���9ن�9ш�9׎�9̗�9l��9h��9\��9B��9O��9.��9��9��9W��9���9��9��9o��9\��9P��9���9���9=��9t��9>y�9�|�9x   x   ,}�9�z�9ry�9��9J��9ۊ�9���9F��9��9���9���9
��9��9���9g��9��9��9���9���9U��9���9���9#��9���9���9��9f��9Kz�9Y|�9�|�9x   x   �{�9ry�9��9��9��9��9ҋ�9��9��9ș�9B��9Ƞ�9@��9*��9]��9Ȣ�9|��9ߡ�9���9���9���9���9Q��9���9���9m��9�9gx�9oz�9�|�9x   x   ��9��9��9���9ˉ�9Ď�9���9���9[��9 ��9Ԝ�9-��9���9���9���9��9��9���9��9W��9��9+��9N��9��9���9{��9��9C��9n~�9O}�9x   x   ���9J��9���9ˉ�9p��9��9k��9i��9��9���9���9��9��9Ҝ�9g��9��9��9l��9��9���9��9���9���9���9���9̃�9���9q��9~��9܃�9x   x   ֆ�9݊�9��9ǎ�9���9&��9���9���9���9��9Ġ�9��9#��9m��9Z��9���9���9;��9���9	��9b��9��9؎�9��9���9���9Ѕ�9ф�9+��9��9x   x   ψ�9���9ϋ�9���9k��9���9���9���9k��9`��9�9@��9 ��9x��9c��9���9���9z��9��9���9*��9��9z��9݉�9���9���9���9֌�9���9��9x   x   Ҏ�9B��9��9���9l��9���9���9���9(��9 ��9��9���9���9���9��9���9��9���9���9��9���93��9|��9H��9X��9��9/��9 ��9��9��9x   x   ͗�9��9��9V��9���9���9k��9#��9V��9]��9M��9w��9���9$��9Y��9o��9<��9+��9���9 ��9��9l��9y��9��9���9N��9���96��9a��9���9x   x   k��9���9Ǚ�9��9���9��9a��9��9a��9U��9��9���9���9h��9���9���9ۘ�9���9̝�9��9H��9<��9��9B��9Q��9��9?��9���9��9���9x   x   d��9���9@��9Ҝ�9���9 �9���9��9J��9��9���9��9ě�9���9Ǜ�9��9	��9R��9���9)��9��9��9��9���9j��9��9���9��9���9���9x   x   [��9��9Ơ�9)��9��9��9D��9���9s��9���9$��9,��9���9���9��9��9���9ǡ�9��9���9X��9���9���9B��9���9p��9���9?��9F��9?��9x   x   B��9ۢ�9A��9 �9��9$��9���9���9���9���9�9���9���9��9â�9}��93��9}��9���9���9���9R��9��9:��9���9q��9{��9S��9���9V��9x   x   Q��9���9+��9���9Ҝ�9i��9y��9���9&��9g��9���9���9��9���9Ť�9��9 ��9���9���9H��9E��9���9���9Ϊ�9���9���9̧�9h��9$��9ͣ�9x   x   +��9k��9]��9���9g��9Y��9d��9��9`��9���9ɛ�9��9¢�9Ƥ�9��9��9��92��9���9��9���9���9ϰ�9!��9��9���9N��9��9W��9���9x   x   ��9��9΢�9��9��9���9���9���9p��9���9��9��9���9��9��9K��97��9o��9���9���9���9���9���98��9l��9��9���9���9��9ߨ�9x   x   ��9��9v��9��9���9���9���9��9<��9ޘ�9��9��9-��9$��9��9:��9���9���9��9���9���9d��9���9 ��9t��9���9!��9���9��9Q��9x   x   Y��9���9ڡ�9���9g��97��9z��9���9*��9���9R��9ǡ�9|��9���9,��9p��9���9Ϯ�9���9���9��9<��9��9ַ�9l��9y��9���9K��9���9���9x   x   ���9���9���9���9��9���9��9�9���9Ν�9���9��9���9���9���9���9��9���9��9d��9Q��9���9��98��9��93��9��9n��9ث�9���9x   x   ��9T��9���9R��9���9��9���9!��9���9��9,��9���9���9M��9��9���9���9���9j��9D��9��9ڻ�9ƺ�9���9���9v��9m��9|��9���9j��9x   x   ��9���9���9��9��9d��9*��9���9��9J��9��9`��9���9E��9���9���9���9��9T��9��9��9��9���9���9��9���9��9��9 ��9��9x   x   p��9���9���9(��9���9��9��95��9l��9?��9	��9���9R��9���9 ��9���9k��97��9ŷ�9ջ�9��9��9µ�9���9$��9��9ʧ�9��9՞�9��9x   x   e��9$��9R��9N��9���9َ�9}��9���9}��9��9��9���9��9���9̰�9���9���9��9��9ź�9���9ȵ�9 ��9ٱ�9(��9G��9w��9��9���9\��9x   x   V��9���9���9���9���9��9��9R��9��9D��9���9G��9:��9̪�9!��9:��9$��9з�9<��9���9���9���9ڱ�9���9ƪ�9X��9��9���9L��9Ő�9x   x   ���9���9���9ʀ�9���9���9���9\��9���9T��9n��9��9��9���9��9k��9z��9k��9��9���9��9 ��9+��9Ǫ�9G��9��9���9���9��9���9x   x   ���9��9n��9|��9̃�9���9Ê�9��9P��9��9	��9r��9n��9���9���9��9���9|��98��9y��9���9��9J��9W��9��9��9���9G��9���9'��9x   x   ;��9l��9ā�9���9���9ԅ�9���9+��9���9@��9���9���9}��9ͧ�9O��9���9��9���9��9k��9��9Ƨ�9x��9��9���9���9���9r��9$��95��9x   x   t��9Jz�9ex�9K��9q��9؄�9֌�9���9;��9���9}��9E��9X��9c��9��9���9���9K��9o��9|��9��9��9��9���9���9J��9s��9��9���9���9x   x   :y�9V|�9kz�9p~�9|��9.��9���9��9c��9��9���9K��9��9*��9[��9	��9��9���9۫�9���9��9ڞ�9���9L��9��9���9%��9���9��9[~�9x   x   �|�9�|�9�|�9Q}�9ك�9��9��9��9���9���9���9E��9T��9Σ�9���9��9Q��9���9 ��9k��9��9��9[��9Ð�9���9(��92��9ۃ�9[~�9�}�9x   x   �I�9�B�9!E�9�G�9�F�9oI�9
M�9<P�9>R�9[�9;Y�9>_�9Ld�9ze�9�g�9c�9�e�9*f�94d�9^�9�Y�96Y�9�R�9&R�9�M�9�I�9 E�9PH�9tB�9�B�9x   x   �B�9�G�9G�9�E�9H�9gN�9ZQ�9�S�9�W�9�Y�9�\�9�]�9/a�9�e�9�d�9�e�9g�9`�9�^�9w\�9W[�9%Y�9�P�9zQ�9|M�9�H�9,F�9�H�94I�9�A�9x   x   $E�9G�9B�9�H�9�I�9�N�9�P�9�V�9�X�9_�9�`�9W^�9e�9b�9r]�9,a�9Vd�9	_�9�`�9�]�9 W�9�W�9�Q�9�N�9.J�9RI�9�?�9�E�92E�9�<�9x   x   �G�9�E�9~H�9�R�9M�9�O�9�R�9zS�9VU�9
Y�9^[�9,_�9�_�9,_�9�_�9f`�9F`�9Y�9�Z�9�W�9�R�9\R�9�N�9|N�9�P�9�I�9BH�9=G�9G�9�F�9x   x   �F�9H�9�I�9M�9�H�9�O�9�U�9�[�9�^�9�^�9^[�9�\�9V_�9�a�9P_�9�[�9\�9`�9�[�9�[�9}V�9�O�9IH�9^M�9�J�9�E�9>F�9�C�9�G�96D�9x   x   iI�9eN�9�N�9�O�9�O�9�R�9�Z�9X�9�[�9�\�9�Y�9^�9�_�9'_�9_�9�Y�9�[�9�\�9�Y�9�Y�9R�9�P�9�N�9O�9�N�9�I�9I�9E�9�D�9�G�9x   x   M�9]Q�9�P�9�R�9�U�9�Z�9KX�9�V�9�[�9�^�9�^�98^�9v\�9A^�9�^�9=_�9�Z�9�V�9
W�9a\�9-T�9�R�9�Q�9�O�9bN�9+N�9�L�9-I�9uM�9oO�9x   x   :P�9�S�9�V�9xS�9�[�9X�9�V�9b�9�`�9�[�9H^�9+a�9ya�9�]�9�[�9�a�9rb�9�V�9X�9�[�9�T�9�U�9JT�9�P�9ER�9	N�9�O�9�O�9�L�9?S�9x   x   3R�9�W�9�X�9QU�9�^�9�[�9�[�9�`�9�Y�9Q^�9�_�9`�9�_�9H_�9xX�9`�9�[�9~]�9 ]�9U�9�X�90W�9lR�9tU�9�T�9�R�9V�9�S�9T�9�U�9x   x   [�9�Y�9_�9Y�9�^�9�\�9�^�9�[�9R^�9[a�9Q]�9�]�9�`�9�^�9c]�9>_�9�Z�9B_�9�[�9�]�9�[�9�Z�9�[�9qX�9�Z�9�T�9�S�9Y\�9X�9�[�9x   x   BY�9�\�9�`�9][�9_[�9�Y�9�^�9H^�9�_�9Q]�9D]�9l]�9�_�9K]�9�\�9V\�9@\�9!Y�9�_�9�\�9�W�9�_�9Y�9�W�9�^�9W�9�]�92W�9fY�9e_�9x   x   :_�9�]�9X^�9+_�9�\�9^�99^�9.a�9#`�9�]�9i]�92`�9Ga�9�`�9^]�9�Z�9�`�98_�9�^�9_�9�_�9|c�9�^�9Nb�9�a�9�c�9�b�9~_�9�c�9�^�9x   x   Gd�91a�9e�9�_�9U_�9�_�9y\�9a�9�_�9�`�9�_�9Fa�9�Z�9�_�9Ca�9�_�9Rd�9�_�9<c�9Vf�9`�91c�9�d�9�d�9�f�9�b�9e�9�a�9�a�9�e�9x   x   ze�9�e�9b�9)_�9�a�9"_�9B^�9�]�9G_�9�^�9K]�9�`�9�_�9W`�9&_�9�a�9g�9g�9
h�99h�9�d�90i�9Ad�9�g�9Oh�9�e�9 j�9xd�9�g�9�g�9x   x   yg�9�d�9n]�9�_�9R_�9_�9�^�9�[�9wX�9_]�9�\�9f]�9Fa�9&_�9�]�9�d�9Qe�9�c�9je�9�j�9�p�9ko�9�n�9�l�9Vn�9m�9|q�9j�9ef�9�d�9x   x   c�9�e�9+a�9c`�9�[�9�Y�9>_�9�a�9	`�9=_�9U\�9�Z�9�_�9�a�9�d�9/d�9Vd�9�j�9h�9�m�9�i�9�j�9Om�9�l�9�l�9wj�9�m�9�h�90i�9c�9x   x   �e�9g�9Xd�9D`�9\�9�[�9�Z�9wb�9�[�9�Z�9C\�9�`�9Qd�9g�9Se�9[d�98k�9�i�9�n�9�k�9l�9�l�97q�9\l�9)k�9(k�9�n�9�i�9�m�9�d�9x   x   )f�9`�9_�9Y�9`�9�\�9�V�9�V�9}]�9?_�9"Y�9=_�9�_�9g�9�c�9�j�9�i�9�r�9�r�9�o�9�s�9zs�9�t�9Us�9%q�9"s�9�r�9&i�9eh�9�d�9x   x   0d�9�^�9�`�9�Z�9�[�9�Y�9W�9X�9]�9�[�9�_�9�^�9<c�9h�9ge�9h�9�n�9�r�9�s�9u�9�v�9�q�97v�9u�9�r�9br�9�o�99i�9Xf�9�g�9x   x   ^�9w\�9�]�9�W�9�[�9�Y�9d\�9�[�9U�9�]�9�\�9_�9Yf�9;h�9�j�9�m�9�k�9�o�9u�9�u�9�u�9qu�9;v�9u�9�q�9Uk�9Wl�9�j�9Sg�9�f�9x   x   �Y�9_[�9W�9�R�9zV�9R�9.T�9�T�9�X�9�[�9�W�9�_�9`�9�d�9�p�9�i�9l�9�s�9�v�9�u�9�z�9pu�9Pv�9&s�9~j�9�k�91q�9�d�9#a�9�_�9x   x   5Y�9#Y�9�W�9aR�9�O�9�P�9�R�9�U�91W�9�Z�9�_�9�c�9.c�91i�9po�9�j�9�l�9�s�9�q�9tu�9xu�9r�9Ot�9�m�9k�9�m�9Fi�9�b�9�b�9X_�9x   x   �R�9�P�9�Q�9�N�9JH�9�N�9�Q�9GT�9kR�9�[�9Y�9�^�9�d�9Fd�9�n�9Jm�97q�9�t�96v�97v�9Mv�9Lt�9�o�96m�9�n�9�e�9�d�9`_�9~Z�9f\�9x   x   #R�9{Q�9�N�9|N�9YM�9O�9�O�9�P�9vU�9vX�9�W�9Kb�9�d�9�g�9�l�9�l�9bl�9Zs�9u�9u�9+s�9�m�9>m�9Ql�9h�9�b�9�b�9�V�9W�9%U�9x   x   �M�9�M�90J�9�P�9�J�9�N�9^N�9BR�9�T�9�Z�9�^�9�a�9g�9Rh�9Xn�9�l�9+k�9%q�9�r�9�q�9�j�9k�9�n�9h�9�f�9|c�9�^�9\�9mV�9XP�9x   x   �I�9�H�9LI�9�I�9�E�9�I�9,N�9N�9�R�9�T�9W�9�c�9�b�9�e�9m�9sj�9*k�9$s�9]r�9Pk�9�k�9�m�9�e�9�b�9~c�9�T�9�T�9~P�9O�9�O�9x   x   E�9,F�9�?�9BH�98F�9 I�9�L�9�O�9V�9�S�9�]�9�b�9
e�9j�9|q�9�m�9�n�9�r�9�o�9Wl�92q�9Gi�9�d�9�b�9�^�9�T�9W�9�O�9K�9[I�9x   x   OH�9�H�9�E�9?G�9�C�9E�9,I�9�O�9�S�9]\�94W�9~_�9�a�9d�9j�9�h�9�i�9$i�9<i�9�j�9�d�9�b�9[_�9�V�9\�9~P�9�O�9YJ�9EE�9UD�9x   x   zB�96I�93E�9�G�9�G�9�D�9uM�9�L�9T�9X�9hY�9�c�9�a�9�g�9df�90i�9�m�9dh�9Zf�9Tg�9&a�9�b�9yZ�9W�9jV�9O�9�J�9HE�9G�9?G�9x   x   �B�9�A�9�<�9�F�94D�9�G�9lO�9<S�9�U�9�[�9g_�9�^�9�e�9�g�9�d�9c�9�d�9�d�9�g�9�f�9�_�9X_�9f\�9&U�9WP�9�O�9XI�9VD�9<G�9?�9x   x   �
�9��9�
�9�9l�9��9$�9��9=�9��9�$�9!�9$�9%�9,&�9-)�9%�9�$�9L$�9s �9�$�9��9�9��9��9��9
�9��9��9j�9x   x   ��9��9�9��9��9��9��9��9��9*�9� �9b�9�"�9�"�9�#�9�$�9�#�9"�9�9 �9�9>�9��9��9x�9�93�9��9��9��9x   x   �
�9�9�92�9��9��9��9~�9��9��9��9��9 "�9�#�9%�9�"�9�!�9��9�9��9��9H�9��9�9��9 �9��98�9R�9��9x   x   �9��9.�9��9E�9��9��9A�9��9��9�"�9�#�9] �9@#�9=$�9� �9�$�9�!�9��9!�92�9�9��9��9��9B�9��9q�9�
�9�	�9x   x   j�9��9��9E�9�9�9��9��9J�9��9�"�9�"�9�!�9�"�9J!�92!�9#�9�9A�9��9�9��9�9��9F�9D�9*�9��9N�9��9x   x   ��9��9��9��9�93�9�9��9��9. �9��9� �9�#�9�"�9T"�9 �9	�9��9b�9�9��9o�9�9��9��9��9��9��9��9�9x   x   $�9��9��9��9��9�9`�9��9��9!�9�!�9��9(!�9��9K �9�!�9�9��9b�9��9��9
�9�9��9��9��92�9^�9�9��9x   x   ��9��9x�9<�9��9��9��9u�9��9!�9�9��9
 �9O�9!�9a�9��9;�9V�9��9>�9��9W�9:�9B�9?�9��9��9��9W�9x   x   ?�9��9��9��9K�9��9��9��9i!�9��9��91�9�9� �9 �9$�98�9��9��9��9=�9��9��9��9'�9�9��9	�9�9�9x   x   ��9"�9��9��9��9. �9!�9!�9��9�!�9f �9]!�9$!�9��9�"�9� �9��9��9��97�9��9��9��9�9��9�9�9��9��9N�9x   x   �$�9� �9��9�"�9�"�9��9�!�9�9��9d �9k�9� �9Y�96�9 �95!�9�"�9�!�9��9o �9$$�9� �9�9k�9�#�9�$�9=#�9��9�9� �9x   x   !�9b�9��9�#�9�"�9� �9��9��9.�9Y!�9} �9�9��9� �9� �9f!�9�$�9 �9��9� �9� �9�#�9��9z�9��9 �9��9� �9d#�9r�9x   x   $�9�"�9"�9[ �9�!�9�#�9&!�9 �9�9)!�9\�9��9S �9@#�9�!�9� �9�!�9�!�9W$�9 �9�#�9-%�9S'�9�'�9<"�9�%�9�&�9�#�9�%�9o �9x   x   %�9�"�9�#�9F#�9�"�9�"�9��9M�9� �9��94�9� �9D#�9�"�9�#�9X#�9\#�9%�9H$�9�(�9S(�9�'�9w*�9�'�9)�9W,�9�(�9�'�9|'�9�#�9x   x   /&�9�#�9%�9?$�9J!�9U"�9K �9!�9 �9�"�9 �9� �9�!�9�#�9!%�9A$�9�%�9E&�9(�9�&�9�%�9+'�97)�9�(�9�'�9�$�9�&�9�&�9�)�9�&�9x   x   ,)�9�$�9�"�9� �9.!�9 �9�!�9e�9*�9� �92!�9`!�9� �9Z#�9A$�9�(�9�*�9<0�9�-�95+�9�/�9�0�9M1�9@1�9�2�9^0�9�*�9.�9�.�9**�9x   x   %�9�#�9�!�9�$�9#�9�9�9��95�9��9�"�9�$�9�!�9]#�9�%�9�*�9�%�9�'�9�-�9C/�9~6�9B1�9�/�9�0�95�9�.�9/.�9r'�92(�9�*�9x   x   �$�9"�9��9�!�9�9��9��9=�9��9��9�!�9 �9�!�9 %�9F&�990�9�'�9�,�9j.�9,�90�9D3�9�3�9�/�9s-�9y.�9�,�9n'�9H.�9 '�9x   x   J$�9�9�9��9B�9c�9c�9V�9��9��9��9��9X$�9I$�9(�9�-�9�-�9m.�9�3�9�1�9�3�9�5�9L3�92�9V2�9.�9R.�9s.�9:)�9D$�9x   x   p �9 �9��9 �9��9�9��9��9��97�9s �9� �9 �9�(�9�&�9:+�9?/�9",�9�1�9�/�9Q1�9q1�9v/�9x1�9/.�9�.�9W*�9'�91'�9[ �9x   x   �$�9
�9��95�9�9��9��9B�99�9��9&$�9� �9�#�9Y(�9�%�9�/�9}6�9
0�9�3�9P1�9D6�9>1�9�3�9�/�9�4�91�9&�9�(�9P%�9� �9x   x   ��9A�9D�9�9��9i�9	�9��9��9��9� �9�#�9.%�9�'�9''�9�0�9C1�9H3�95�9u1�9C1�9Z5�9h3�9�1�9�1�9&�9g'�9�$�9:"�9� �9x   x   �9��9��9��9
�9!�9�9[�9��9��9�9��9W'�9t*�99)�9M1�9�/�9�3�9K3�9r/�9�3�9g3�9&/�9+1�9	(�9�+�9�'�9< �9� �9��9x   x   ��9��9�9��9��9��9��9>�9��9�9j�9~�9�'�9�'�9�(�9D1�9�0�9�/�9 2�9y1�9�/�9�1�9.1�9)�9�(�9�%�9��94�9��9I�9x   x   ��9y�9��9��9F�9��9��9H�9(�9��9�#�9��9?"�9)�9�'�9�2�95�9r-�9X2�9-.�9�4�9�1�9(�9�(�9�!�9l�9�#�9��9�9{�9x   x   ��9�9"�9G�9C�9��9��9@�9�9 �9�$�9�9�%�9U,�9�$�9g0�9�.�9�.�9.�9�.�91�9!&�9�+�9�%�9n�9F"�9��9��9��9a�9x   x   �93�9��9��9,�9��94�9��9��9	�9=#�9��9�&�9(�9�&�9�*�9/.�9�,�9X.�9U*�9&�9h'�9�'�9��9�#�9��9��9�9"�9��9x   x   ��9��97�9r�9��9��9\�9��9�9��9��9� �9�#�9�'�9�&�9 .�9p'�9j'�9o.�9'�9�(�9�$�9@ �96�9��9��9	�9�9��9��9x   x   ��9��9R�9�
�9S�9��9�9��9�9��9�9a#�9�%�9y'�9�)�9�.�92(�9M.�98)�91'�9M%�9;"�9� �9��9�9��9$�9��9��9I
�9x   x   c�9��9��9�	�9��9!�9��9]�9�9J�9� �9t�9p �9�#�9�&�9(*�9�*�9'�9E$�9\ �9� �9� �9��9J�9y�9d�9��9��9J
�9��9x   x   ���9z��9���9��9���9N��9���9���9���9���9���9���9j��9���9���9���9���9}��9���9t��9���9���9���9��9N��9
��9Q��9{��9���9^��9x   x   y��9���9���9���9���9���9���9E��9���9���9���9P��9���9���9���9��9���9���9d��9���9_��9���9l��9���9*��9q��92��9���9���9���9x   x   ���9���9T��9��9p��9C��9<��9���9���9_��9[��9���9���9��9��9��9��9:��9n��9(��9���9��9���9y��9���9���9*��9w��9���9$��9x   x   ��9���9	��9~��9}��9���9���9���9���9���9��9��9��9���9���9;��9���9���9o��9���9B��9���9!��9���9���96��9���9U��9y��9-��9x   x   ���9���9p��9x��9*��9G��9��9���9��9���9���9���9���9{��9Z��9+��94��9���9I��9���9n��9���9
��9���9���9q��9���9��9H��9���9x   x   O��9���9F��9���9A��9c��9[��9���9���9���9!��9D��9��9q��9M��9!��9���9���9&��9���9���9���9��9��9���9���9o��9���9]��9���9x   x   ���9���9;��9���9��9_��9c��9���9���9E��9���9���9���9���9���9��9���9���9V��9&��9^��98��9���9���9���9���97��9���9���9���9x   x   ���9A��9���9���9���9���9���9y��9c��9o��9���9{��9���9���9���9��9���9��9=��9P��9��9U��9��9d��9���9���9���9��9���9&��9x   x   ���9���9���9���9��9���9���9g��9���9���91��9���9��9i��9L��90��9���9���9���9���9��9���9��9#��9t��9���9���9���9l��9���9x   x   ���9���9`��9���9���9���9@��9q��9���9���9��9s��97��9)��9���9���9���9/��9K��99��9���98��9���9���9#��9���9��9D��9��9��9x   x   ���9���9^��9��9���9 ��9���9���93��9��9���9/��9��9t��9"��9y��9���9%��9���9���9���9%��9���9Y��9'��9���9���9���9���9{��9x   x   ���9M��9���9��9���9F��9���9���9���9y��90��9��9p��9���9���9���9]��9l��9���9h��9o��9���9W��9���9���9���9���9���9���9���9x   x   m��9��9���9 ��9���9��9���9���9��94��9��9p��9��9y��9+��9G��9���9���9��9���9}��9u��9��9q��9j��9��92��9���9���9R��9x   x   ���9���9��9���9s��9m��9���9���9e��9'��9u��9���9x��9>��9��9���9���9���9^��9���9H��9���9 ��9���9H��9���9���9���9+��91��9x   x   ���9���9
��9���9W��9K��9���9���9H��9���9$��9���9*��9��9���9,��9o��9���9���9;��9l��9���93��9��9���9%��9���9Z��9��9���9x   x   ���9��9��9A��90��9%��9��9��9,��9���9���9���9L��9���90��9��9��9���9
��9^��9���93��9���9���9E��9��9���9#��9���9��9x   x   ���9���9��9���95��9���9���9���9���9���9���9^��9���9���9s��9��9���9���9���9���9o��9��9���9���9n��9���9d��93��9���9���9x   x   ~��9���93��9���9���9���9���9��9���9,��9$��9g��9���9���9���9���9���9���9��9���9>��9l��9��9���9��9���9���9���9x��9C��9x   x    ��9a��9r��9o��9E��9+��9V��9?��9���9L��9���9���9��9_��9���9��9���9��9���9:��9;��9_��9V��9h��97��9���9��9��9���9���9x   x   y��9���9-��9���9���9���9#��9T��9���9=��9���9h��9���9���9:��9[��9���9���9<��9)��9��9���9o��9���9���9���9��9i��9���9���9x   x   ���9Y��9���9B��9o��9���9_��9��9��9���9���9s��9|��9F��9n��9���9s��9?��9<��9��9���9 ��9<��9��9e��9���9b��9���9H��9*��9x   x   ���9���9��9���9���9���97��9T��9���92��9%��9���9w��9���9���93��9��9h��9_��9}��9���9-��9���9{��9���9��9���9���9$��9���9x   x   ���9i��9���9!��9��9��9���9��9��9���9���9V��9��9%��95��9���9���9��9[��9r��9?��9���9B��9���9 ��9���9���9���9���9���9x   x   ��9���9}��9���9���9��9���9c��9'��9���9b��9���9o��9���9��9���9���9���9h��9���9��9z��9���9���9L��9���9w��9���9$��9���9x   x   O��9(��9���9���9���9���9���9���9v��9%��9(��9���9m��9M��9���9D��9r��9��98��9���9e��9���9"��9O��9g��9��9���9q��9Z��9���9x   x   	��9p��9���94��9r��9���9���9���9���9���9���9���9��9���9&��9��9���9���9���9���9���9��9���9���9��9
��9���90��9A��9$��9x   x   R��93��9'��9���9���9p��9>��9���9���9��9���9���94��9���9���9���9_��9���9���9��9a��9���9���9t��9���9���93��9���9���91��9x   x   |��9���9w��9V��9��9���9���9��9���9F��9���9���9���9���9_��9'��98��9���9��9p��9���9���9���9���9o��9/��9���9���9���9��9x   x   ���9���9���9z��9H��9X��9���9~��9k��9	��9���9���9���9/��9��9���9���9v��9���9���9K��9%��9���9#��9X��9A��9���9���9���9 ��9x   x   ]��9���9#��9,��9���9���9���9%��9���9��9z��9���9R��95��9���9
��9���9A��9���9���9)��9���9���9���9���9"��9.��9��9���9���9x   x   3��9ϗ�9q��9���9ٙ�9���9���9���9J��9w��9��9��9+��9��9^��9���9-��9Ʃ�9z��9G��9D��9���9���9���9*��9��9`��9���9��9��9x   x   җ�9���9���9���9
��9���9e��9���9���9���9���9'��9���98��9��9i��96��9���9���9?��9��9��9Ǡ�9���9z��9Q��9��9���9���9��9x   x   t��9���9��9���9���9���9Ȥ�9���9���9!��9���9:��9Y��9ƨ�9t��9���9m��9k��9���9��9��9���9r��9A��9��9ʜ�9~��9G��9Җ�9^��9x   x   ���9���9��9Q��9��9���9��9��9{��9.��9���9��9ت�9��9z��9���9��9x��9Ϣ�9���9l��9��9r��9&��9���96��9;��9���9~��9���9x   x   ڙ�9	��9���9��9��9N��9���9��96��9���9��9��9��9$��9���9���9'��9/��9���9*��9��9ȡ�9���9��9���9��9�9C��9Ϡ�9{��9x   x   ���9���9���9���9N��9��9���9���9��9��9`��90��9ϫ�9��9#��9���92��9ƥ�9_��9��9��9���9��9-��9d��9؜�9���9ƛ�9]��9��9x   x   ���9h��9Ȥ�9��9���9���9*��9���9���9ר�9n��9H��9���9���9Ũ�9"��9Ш�9ˡ�9G��9ߤ�9��9���9��9B��9��9���9ڡ�9��9���9���9x   x   ��9���9���9��9��9���9���9M��9l��9ѥ�9���9Ʀ�96��9	��9ץ�9���9���9���9J��9���9��9���9���92��9}��9K��9N��9���9d��9ȟ�9x   x   G��9���9���9|��98��9	��9���9o��9ĥ�9r��9���9���9���9i��9I��9���9`��9���9���9v��9���9ߢ�9[��9���9S��9o��9ӡ�9ͣ�9.��9У�9x   x   s��9���9��9.��9���9��9ب�9ҥ�9o��9��9��9���9~��9��9���9���9��9���9��9S��9$��9���9#��9٣�9 ��9��9A��9���9K��9\��9x   x   ��9���9���9���9��9c��9p��9���9���9��9���9��9���9���9��9y��9ʩ�9��9J��91��9���9Ӭ�9���9k��9��94��9���9���9���9b��9x   x   ��9%��96��9��9��90��9D��9Ŧ�9���9���9��9B��9L��9���9���9���9��9M��9G��9=��9ܬ�9���9��9��9��9 ��9q��9���9-��9���9x   x   *��9���9Z��9ת�9��9Ϋ�9���95��9���9��9���9M��9���9���9���9���9���9���9���9S��9���9Ϋ�9���9ө�9D��9)��9[��9N��9��9|��9x   x   ���96��9¨�9��9-��9��9���9
��9l��9��9���9���9���9���9*��9���9���9(��9���9ʨ�9���9Ѯ�9Z��9���9���9��9U��9U��9~��9���9x   x   ]��9��9r��9~��9���9%��9Ĩ�9ץ�9M��9���9��9���9���9,��96��9���9��9#��9��9���9���9���9���9���9��9���9��9���9��9���9x   x   ���9h��9���9���9y��9���9!��9���9���9���9y��9���9���9���9���9���9d��9��9j��9f��9��9��9���9���9���9ˮ�9���9l��9O��9��9x   x   '��95��9p��9���9#��94��9Ԩ�9���9f��9��9ũ�9��9���9���9��9h��9���9Ӯ�9\��90��9��9��9��9��9���9q��9%��9���9)��9I��9x   x   ĩ�9���9o��9z��91��9ĥ�9ˡ�9���9���9ħ�9	��9T��9§�9(��9 ��9��9ծ�9/��9���9���9^��9��9V��9��9˳�9���9���9r��9"��9���9x   x   y��9���9���9Ϣ�9���9\��9I��9H��9���9��9M��9F��9���9���9��9c��9a��9���9���9��9޴�9`��9��9���9���9r��9���9��9��9��9x   x   @��9;��9��9���9,��9��9��9���9u��9R��9-��9<��9S��9Ҩ�9���9j��97��9���9��96��9ȴ�9��9��9���9���9���9��9İ�9$��9A��9x   x   H��9��9��9j��9��9��9��9��9���9(��9���9ެ�9���9���9���9��9��9_��9޴�9̴�9��9ʹ�9��9���9���9��9��9%��9��9��9x   x   ���9��9���9��9ȡ�9���9���9���9��9���9Ь�9��9Ы�9Ю�9���9ݱ�9��9��9_��9��9˴�9|��9���9ݵ�9G��9̴�9s��9���9���9#��9x   x   ���9Ơ�9v��9r��9���9���9��9���9a��9'��9���9��9���9\��9���9���9���9X��9��9��9��9���9ĵ�9��9��9���9��9"��9��9q��9x   x   ���9���9B��9%��9��9.��9C��9.��9���9գ�9j��9��9Щ�9���9���9���9��9��9���9���9���9��9��9���9#��9}��9���9o��9��9գ�9x   x   ,��9~��9��9���9���9g��9��9z��9T��9���9	��9��9E��9���9��9���9���9˳�9���9���9���9M��9��9#��9���97��9q��9���9w��9���9x   x   "��9T��9˜�95��9��9ۜ�9���9K��9v��9��9:��9$��9%��9��9���9Ů�9w��9���9s��9���9��9ʹ�9���9~��98��9���9���9פ�9���91��9x   x   ]��9��9���9;��9���9���9ء�9I��9ա�9<��9���9v��9X��9W��9��9���9,��9���9���9��9!��9v��9��9ì�9o��9���9��9Y��9��9���9x   x   ���9���9K��9���9?��9Ǜ�9��9��9ң�9���9���9���9M��9R��9���9g��9���9v��9��9���9%��9���9!��9t��9���9դ�9_��9��9U��9���9x   x   ��9���9і�9���9Ҡ�9`��9���9d��9-��9K��9���91��9��9}��9	��9O��9'��9!��9��9��9��9���9��9���9w��9���9��9X��9��9\��9x   x   ��9��9]��9���9��9��9���9ɟ�9ϣ�9_��9a��9���9}��9���9~��9��9F��9���9��9B��9��9%��9q��9ԣ�9���92��9���9���9\��9_��9x   x   %c�9�c�9?b�9�_�9:f�9�g�9�d�9Ok�9�k�9hi�9�k�9�p�9rs�94q�9�m�9�o�9�n�9�p�9s�9q�93l�9�j�9!k�9j�92d�9�g�9g�9_�9�d�9�c�9x   x   �c�9~_�9+c�9f�9�e�9�c�9�f�9Ok�9jm�9~j�9Br�9�r�9�o�9p�9r�9Pq�9�n�9'q�9�q�9_r�9Xi�9Ml�9[m�9g�9 d�9pe�9pf�9�a�9�]�9Sd�9x   x   <b�9+c�9(d�9�b�9Qf�97g�9Kh�9�i�9�l�9Hl�9�o�9�n�9Ol�9�m�9v�9�n�9rl�97n�9�o�9�l�9n�9[i�9�f�9�g�9�f�9�a�9�e�9!d�9�b�9�i�9x   x   �_�9 f�9�b�9Jb�9c�9�e�9�e�9?n�9Co�9m�9En�98p�9�n�9�r�9�q�9=n�9ho�9�o�9gl�9*n�9(n�9�e�9�f�9�a�9�c�9�a�9�d�9�_�9�`�9b�9x   x   <f�9�e�9Sf�9
c�9�j�9�j�9Gh�9�l�9k�9`m�9<o�9�k�9sm�9Hl�9lm�9jm�9o�9l�9m�9�l�9^h�9�j�9k�9yb�9f�9�g�9.f�9�^�9Pa�9E^�9x   x   �g�9�c�94g�9�e�9k�9ph�9�f�9�m�9dj�9Yk�90m�9:p�9~k�9zl�9�n�95l�9�l�9-j�9�l�91g�9h�9�i�98g�9�f�9Lc�9 g�9�g�9�e�9�e�9oh�9x   x   �d�9�f�9Fh�9�e�9Fh�9�f�9�m�9Aq�9�j�9�l�9�n�9�n�9|m�9�n�9Ip�9{l�9�j�9pq�9�n�9�e�9ej�9�d�96g�9Ch�9�c�98f�9�c�9Qb�9Yd�9�d�9x   x   Kk�9Ok�9�i�9@n�9�l�9�m�9Dq�9j�9Uj�9�p�9�k�9jp�9xo�9fk�9�p�9�i�98j�9\q�9�m�9l�9Tm�9�j�9k�9k�9�i�9�e�9�j�9;j�9�f�9�i�9x   x   �k�9km�9�l�9Fo�9k�9dj�9�j�9Pj�9�m�9�n�9`l�9Uo�9�m�9�m�9�n�9�j�9Fj�9�i�9�l�9Ko�9m�9~m�9�k�9`l�9Fh�9vf�9�k�9�e�9�h�9�k�9x   x   di�9�j�9Gl�9m�9]m�9Yk�9�l�9�p�9�n�9�n�9?o�9n�9�n�9(o�9�n�9�l�9�l�9*l�9�k�9�l�9i�9
j�9�j�9�i�9k�9�g�93i�9j�9�i�9�j�9x   x   �k�9Dr�9�o�9In�9=o�90m�9�n�9�k�9el�9>o�9�u�9+o�9;l�9�l�9�p�9vk�9 o�9�o�9 p�9~r�9�l�9�p�9�o�9�m�9�p�9Ol�9�p�9�n�9�o�9Fq�9x   x   �p�9�r�9�n�9=p�9�k�97p�9�n�9hp�9Zo�9
n�9)o�9�o�9�o�9Tm�9#p�9m�9�o�9n�9r�9�p�9�i�9l�9}m�9el�9�l�93k�9Kl�9�l�9l�9Jk�9x   x   rs�9�o�9Ll�9�n�9pm�9|k�9m�9vo�9�m�9�n�9<l�9�o�9o�9�k�9]m�9n�9�l�9�p�9�s�9�r�9vq�9At�9�s�9Mq�9Ao�9cs�9(s�9�u�9p�9�q�9x   x   /q�9p�9�m�9�r�9@l�9vl�9�n�9ck�9�m�9#o�9�l�9Pm�9�k�9Ml�9Wr�9�n�9o�9vp�9Uo�97r�9}u�9�p�9�s�9�w�9)v�9�r�9p�9Wu�9�s�9�o�9x   x   �m�9r�9v�9�q�9hm�9�n�9Jp�9�p�9�n�9�n�9�p�9#p�9\m�9Zr�9�u�9�q�9�n�9`o�9s�9�r�9|n�9�m�9�o�96u�9�p�9'p�9�m�9�r�9�q�9�n�9x   x   �o�9Pq�9�n�9>n�9lm�95l�9}l�9�i�9�j�9�l�9xk�9m�9n�9�n�9�q�9�o�9�r�9�t�9|w�9br�9�x�9�y�9�s�9�t�9jw�9�w�9�s�9%w�9�u�9�s�9x   x   �n�9�n�9ol�9po�9o�9�l�9�j�90j�9Fj�9�l�9!o�9�o�9�l�9o�9�n�9�r�95t�9r�9zv�9'w�9�w�9�v�9 r�9.w�9�y�9Bw�9�u�9�r�9�q�9�r�9x   x   �p�9 q�92n�9�o�9l�9+j�9rq�9Xq�9�i�9/l�9�o�9n�9�p�9yp�9do�9�t�9r�9�s�9Uu�9�v�9u�9$s�9Cr�9�t�9Au�9Ou�9Yt�9Os�9jv�9�n�9x   x   s�9r�9�o�9dl�9m�9�l�9�n�9�m�9�l�9�k�9p�9 r�9�s�9Uo�9s�9w�9tv�9Ou�9�q�9�z�9�u�9�z�9�v�9+z�9Js�9�u�9u�9�v�9�q�9�o�9x   x   q�9cr�9�l�9,n�9�l�90g�9�e�9l�9Lo�9�l�9�r�9�p�9�r�97r�9�r�9ar�9$w�9�v�9�z�9~v�9�y�9�x�9wv�97{�9<t�9�w�9�s�9Ms�9Bs�9Yr�9x   x   3l�9Xi�9n�9'n�9`h�9h�9ej�9Sm�9m�9	i�9�l�9�i�9wq�9~u�9}n�9�x�9�w�9u�9�u�9�y�9�|�9�y�9)u�9�u�9�y�9+w�9wm�9;u�9 p�9�j�9x   x   �j�9Ll�9Yi�9�e�9�j�9�i�9�d�9�j�9{m�9j�9�p�9}l�9Dt�9�p�9�m�9�y�9�v�9's�9�z�9�x�9�y�9H{�9�r�9v�9�x�9�o�9q�9*u�93m�9Vp�9x   x   !k�9Ym�9�f�9�f�9k�97g�95g�9k�9�k�9�j�9�o�9zm�9�s�9�s�9�o�9�s�9r�9Fr�9�v�9uv�9)u�9�r�9�r�9Tt�9_p�9�r�9�r�9�l�9Yo�9�j�9x   x   #j�9g�9�g�9�a�9~b�9�f�9Gh�9k�9`l�9�i�9�m�9kl�9Xq�9�w�97u�9�t�9)w�9�t�9/z�97{�9�u�9v�9Qt�9;u�9�v�9Cs�9�l�9^n�9qj�9.l�9x   x   /d�9d�9�f�9�c�9f�9Gc�9�c�9�i�9Jh�9k�9�p�9�l�9@o�9)v�9�p�9qw�9�y�9Cu�9Os�9:t�9�y�9�x�9^p�9�v�9[o�9k�9�p�9
j�9g�9�k�9x   x   �g�9le�9�a�9�a�9�g�9g�97f�9f�9sf�9�g�9Pl�9-k�9ls�9�r�9(p�9�w�9<w�9Iu�9�u�9�w�9,w�9�o�9�r�9Bs�9k�9�m�9�g�9?h�9e�9�d�9x   x   g�9mf�9�e�9�d�91f�9�g�9�c�9�j�9�k�96i�9�p�9Ml�9+s�9p�9�m�9�s�9�u�9]t�9u�9�s�9xm�9q�9�r�9�l�9�p�9�g�9Vj�9]j�9ne�9�g�9x   x   _�9�a�9$d�9�_�9�^�9�e�9Pb�9?j�9�e�9j�9�n�9�l�9�u�9Wu�9�r�9$w�9�r�9Ks�9�v�9Ks�9:u�9+u�9�l�9_n�9
j�9Bh�9`j�9�a�9Ce�9.^�9x   x   �d�9�]�9�b�9�`�9La�9�e�9Td�9�f�9�h�9�i�9�o�9l�9p�9�s�9r�9�u�9�q�9qv�9�q�9Js�9#p�97m�9Xo�9pj�9g�9�d�9ie�9>e�9�b�96a�9x   x   �c�9Ud�9�i�9b�9F^�9oh�9�d�9�i�9�k�9�j�9Fq�9?k�9�q�9�o�9�n�9�s�9�r�9�n�9�o�9Vr�9�j�9Yp�9�j�9.l�9�k�9�d�9�g�9*^�96a�9h�9x   x   @,�9(�9q+�9�/�9�-�9=.�9�2�9�.�94�9�4�9U9�9 4�9g5�9�:�9�8�9�;�9c:�9!;�9~4�9�4�9�8�9e6�9�3�9�,�9L3�9�.�9/-�9�.�9�.�9](�9x   x   (�9�-�9�,�9+�9�*�9�0�9�-�9{.�9�4�9�2�9o2�9�0�9:8�9V9�9?6�9�5�9-7�99�9�0�9x2�9�2�9^3�9m0�9q-�9�0�9�*�9,�9�+�9�*�9�'�9x   x   q+�9�,�90-�9Q.�9�0�9�2�951�9`0�9E/�9>0�974�9�5�9]7�9@6�9`4�98�9"8�9�5�9�3�9�0�9 0�9c/�9�0�9�3�9P0�9k-�9�-�9�-�9�-�9�(�9x   x   �/�9+�9Q.�92�9�1�9�3�9�3�9%2�9�3�98�93�9�4�99�96�9�4�9C8�9|3�9)4�9_8�9Q2�9L3�9�3�9Y3�9�0�9�3�9�-�9U*�9�.�9�,�9/�9x   x   �-�9�*�9�0�9�1�9l,�9Q-�9�3�9�0�952�9�5�9�2�9�6�9k6�9�4�9(7�9Z8�93�9�3�9�3�9�0�9�2�9�-�9�,�9�0�9�/�9,�9�-�9F/�9u-�9.�9x   x   8.�9�0�93�9�3�9O-�9�5�9�6�9v1�9�5�9�7�9�5�9K:�907�9<8�9A8�9�4�9m9�905�9�0�9�7�9�5�9T,�9p4�93�9v0�9-�9�+�9-2�9N1�9U,�9x   x    3�9�-�9;1�9�3�9�3�9�6�991�9 2�9e8�9�4�91�9�5�9�5�9�5�9�3�9�3�9�8�9K2�9b1�946�9�4�983�9m0�9/�93�9Z/�9.�9i*�9�/�9�-�9x   x   �.�9y.�9c0�9&2�9�0�9v1�92�9�4�9p8�98�9T5�9�6�9c6�9a4�9�7�918�9�4�9p2�9�1�9t0�9�1�9�1�9�-�9�-�9�/�97�9�1�9e0�9�6�9�/�9x   x    4�9�4�9B/�9�3�962�9�5�9e8�9u8�9�3�9�4�9�6�9g5�9w8�93�9@5�99�98�9�4�9N3�9�3�9�.�9a4�95�9T1�9�0�9�2�9�2�9�2�962�9�/�9x   x   �4�9�2�9:0�98�9�5�9�7�9�4�98�9�4�9f5�9�3�9�1�9m6�9>5�9u5�95�9:9�9�4�9�6�9d1�9w2�95�9n1�9�4�9�2�9&4�9�5�91�9�4�93�9x   x   R9�9k2�994�93�9�2�9�5�91�9Q5�9�6�9�3�9c5�9n3�9c5�9m6�9i3�9�3�9{2�9�4�9�3�9!2�9-:�9�1�937�96�9�4�9�7�9�4�9}7�9�6�9o1�9x   x    4�9�0�9�5�9�4�9�6�9J:�96�9�6�9f5�9�1�9m3�9J6�9�6�94�9�9�9u8�9�3�9p5�9�0�9�3�9f5�9�4�9<:�9�3�9�9�918�9�3�9:�9�3�9�6�9x   x   f5�9:8�9Z7�99�9p6�937�9�5�9b6�9u8�9n6�9f5�9�6�9�6�98�96�9�8�9+8�9�8�9[5�98�9�9�9�2�95�9'7�9�8�9�8�9�3�9�4�9	9�9E7�9x   x   �:�9Y9�9E6�96�9�4�9<8�9�5�9e4�93�9=5�9r6�94�9 8�9�4�9�5�97�98�9:�9Y6�9�7�9�:�9�7�9�=�9`7�9�6�9o=�927�9�9�9�8�9u6�9x   x   �8�996�9a4�9�4�9,7�9@8�9�3�9�7�9?5�9t5�9l3�9�9�96�9�5�9V4�9�5�9B:�9�;�9�7�98�9�?�9�<�9�8�93:�9J8�9�>�9�?�9[8�9+7�9A;�9x   x   �;�9�5�98�9C8�9X8�9�4�9�3�938�99�9�4�9�3�9w8�9�8�97�9�5�9�;�9�8�9�8�9�9�9v8�9=�9#9�9�>�9t@�9H7�9�;�9�9�9�8�9`9�9Z:�9x   x   b:�9/7�9$8�9}3�93�9k9�9�8�9�4�98�979�9{2�9�3�908�98�9E:�9�8�9�5�9�<�9�;�9"9�9A8�9�;�9�>�9=<�9%:�9<9�9;�9�=�93�9�8�9x   x   ;�99�9�5�9(4�9�3�935�9O2�9v2�9�4�9�4�9�4�9q5�9�8�9:�9�;�9�8�9�<�9v=�9�<�9�>�9,=�9�B�9�@�9�<�9�=�9u<�99=�9T=�9�:�9�:�9x   x   ~4�9�0�9�3�9_8�9�3�9�0�9^1�9�1�9K3�9�6�9�3�91�9]5�9W6�9�7�9�9�9�;�9�<�9>�9S?�9�=�9�@�9�?�9�>�9=?�9�=�9�:�9r8�9�6�9�6�9x   x   �4�9r2�9�0�9R2�9�0�9�7�9-6�9s0�9�3�9h1�9 2�9�3�98�9�7�9�7�9u8�9%9�9�>�9S?�9O?�9�<�9�;�9->�9�?�9e<�9M9�9I:�9r8�9�8�9w7�9x   x   �8�9�2�9#0�9K3�9�2�9�5�9�4�9�1�9�.�9u2�9+:�9f5�9�9�9�:�9�?�9=�9?8�9(=�9�=�9�<�9!>�9�<�9<>�9>�9J:�9J;�9?�9�9�9�8�9�6�9x   x   j6�9a3�9h/�9�3�9�-�9U,�9:3�9�1�9d4�95�9�1�9�4�9�2�9�7�9�<�9"9�9�;�9�B�9�@�9�;�9�<�9�@�9�@�9f:�9�8�9,>�9^8�9W4�9�4�9�0�9x   x   �3�9n0�9�0�9Z3�9�,�9p4�9m0�9�-�95�9j1�947�98:�95�9�=�9�8�9�>�9�>�9�@�9�?�9,>�9@>�9�@�9�A�9�>�99�9;<�94�9G9�9�6�92�9x   x   �,�9v-�9�3�9�0�9�0�93�9	/�9�-�9T1�9�4�9�6�9�3�9%7�9c7�97:�9t@�9<<�9�<�9�>�9�?�9>�9g:�9�>�9p:�9
7�99�9�3�9�7�9(5�9�0�9x   x   K3�9�0�9U0�9�3�9�/�9{0�93�9�/�9�0�9�2�9�4�9�9�9�8�9�6�9K8�9H7�9$:�9�=�9@?�9d<�9I:�9�8�99�97�9@8�9|8�9K4�9^1�9F0�9I2�9x   x   �.�9�*�9n-�9�-�9,�9-�9Z/�97�9�2�9)4�9�7�988�9�8�9o=�9�>�9�;�9>9�9t<�9�=�9N9�9K;�9(>�9=<�99�9�8�99�9�4�9K5�95�9�,�9x   x   /-�9,�9�-�9R*�9�-�9�+�9.�9�1�9�2�9�5�9�4�9�3�9�3�977�9�?�9�9�9";�9>=�9�:�9L:�9
?�9_8�94�9�3�9R4�9�4�91�9�0�9b1�9�+�9x   x   �.�9�+�9�-�9�.�9E/�9+2�9k*�9j0�9�2�91�9~7�9:�9�4�9�9�9Y8�9�8�9�=�9Z=�9p8�9r8�9�9�9T4�9H9�9�7�9_1�9K5�9�0�9D)�9�0�9/�9x   x   �.�9�*�9�-�9�,�9y-�9P1�9�/�9�6�922�9�4�9�6�9�3�99�9�8�9*7�9c9�93�9�:�9�6�9�8�9�8�9�4�9�6�9%5�9F0�9	5�9f1�9�0�9�.�9*-�9x   x   `(�9�'�9�(�9/�9.�9Z,�9�-�9�/�9�/�93�9q1�9�6�9H7�9s6�9:;�9U:�9�8�9�:�9�6�9v7�9�6�9�0�92�9�0�9G2�9�,�9,�9/�9,-�9'�9x   x   X��9L��9���9���9���9O��9���9���9���9y��9���9{��9� �9P��9���9 �9���9s��9���9{��9g��9J��9���9��9���9J��9��9��9���9y��9x   x   L��9]��9���9��9h��9Y��9N��9���9E��9z �9���9��98��9���9��9�9���9D��9O�9���9� �9.��9��9Q��9c��9���9���92��9���9F��9x   x   ���9���9&��9���9z��9���9��9���9� �9� �9���9�9h��9[�9��9�9���9��9q��9?�9F�9;��9���9���9a��9���9Z��9C��9	��9���9x   x   ���9��9���9��9i��9���9H��9��9���9��9��9� �9���9R��9���9���9g��9h��9���9p��9���9���9r��94��9���9���9e��9��9���9��9x   x   ���9l��9x��9f��9��9W��9;��9}��9���9���9���9W��9���9\�9���9���9���9��9[��9��9���9���9��9K��9 ��9&��9 ��9���9���9���9x   x   O��9W��9���9���9Y��9���9���95�9/��9���9� �9���9���9s��9F��9 �9*��9O��9� �9���96��9���9Q��9��9���9���9t��9,��9���9���9x   x   ���9I��9��9G��9;��9���9A��9!��9���9���9���9���9���9h��9���9k��9���97��9���9"��9!��9s��9(��9e��9?��9���9O��9���9���9&��9x   x   ���9���9���9��9y��93�9"��9���9��9:��97 �9%��9���9���9c��9���9��9���9b�9���9���9���9���9k��9P��9���9 ��9{��9���9���9x   x   ���9C��9� �9���9���9,��9���9"��9/��9f��9���9���9 �9���9���9���9O��9���9���9���9���9+��9Q��9n��9$��9g��9���9���9���9���9x   x   z��9z �9� �9��9���9���9���99��9c��94��9� �9��9�9���9��93��9���9���9��9��9� �9S��9F��9��9 �9���9���9���9���9m��9x   x   ���9���9���9��9���9� �9���99 �9���9� �9L �9R �9���9b�9R��9+��9��9���9?��9���9���9U��9���9���9���9���9���9���9���9���9x   x   ~��9��9�9� �9W��9���9���9*��9���9��9S �9P��9���9@��9���9{��9��9��9��9��91�9x�9��9��9m �9P��9��9��9��9��9x   x   � �9=��9g��9���9���9���9���9���9 �9�9���9���9���9���9W��9���9���9<��9 �98��9���9u��9��9���9W �9O��9� �9� �92��9S��9x   x   O��9���9X�9N��9]�9q��9f��9���9���9���9a�9A��9���9��9��9n�9���9l��9��9���9M��9� �9� �9T��9���9 �9D �9���97��9?�9x   x   ���9��9��9���9���9H��9���9`��9���9��9P��9���9Z��9!��9
��9��95��9��9��95�9T�9�9��9t�9��9��9=�9�9��9��9x   x    �9�9�9���9���9 �9h��9���9���94��9-��9y��9���9n�9��9���9� �9���9��9��9Q �9q�9R�9y�9�9���9��9l �9& �9��9x   x   ���9���9���9c��9���9*��9���9��9N��9���9��9��9���9���94��9� �9"�9E�9��9��9��9��9K��9�9��9]�9��9��99�9���9x   x   n��9L��9��9n��9��9N��91��9���9���9���9���9��9B��9g��9��9���9C�9���9��9�9��9��9s�9��9��90�9;��9{�9Z�9� �9x   x   ���9N�9n��9���9Y��9� �9���9h�9���9��9<��9��9	 �9��9��9��9��9��9��9l��91�9���9#�9S��9f�9�92�9 �9�9��9x   x   z��9���9?�9n��9��9���9$��9���9���9��9���9��99��9���9:�9��9��9�9j��9��95�9N�9��9n��9��9;�9�9F�9U �9���9x   x   m��9� �9C�9���9���98��9"��9���9���9� �9���92�9���9L��9U�9R �9��9��95�95�9��95�9
�9��9h�9���9v�9���9���9�9x   x   K��9+��98��9���9���9���9r��9���9*��9S��9T��9z�9u��9� �9�9q�9��9��9���9M�90�9��9K�9�9�9��9� �9h �9��9\��9x   x   ���9��9���9s��9��9N��9)��9���9T��9G��9���9��9��9� �9��9Q�9O��9o�9%�9��9
�9E�9]�9 �9��9 �9l�9 �9���9���9x   x   ��9O��9���93��9P��9��9b��9k��9v��9���9���9��9���9W��9p�9w�9�9��9Q��9m��9��9�9�9��9���9���9[�9��9���9 ��9x   x   ���9]��9b��9���9��9���9A��9U��9&��9 �9���9t �9V �9���9��9�9��9��9j�9��9e�9�9��9���9���9���9���9���9���9���9x   x   P��9���9~��9���9"��9���9���9���9n��9���9���9T��9G��9#�9��9���9a�9.�9�9@�9���9��9 �9���9���9���9i��9l��9V��9���9x   x   ��9���9Z��9i��9 ��9t��9Q��9��9���9���9���9��9� �9G �9A�9��9��96��9.�9�9z�9� �9l�9Z�9���9f��9���9���9��9>��9x   x   ���91��9B��9��9���9.��9���9u��9 ��9���9���9��9 �9���9�9h �9��9��9 �9G�9���9h �9 �9��9���9i��9���9T��9���9���9x   x   ���9���9��9���9���9���9���9���9���9���9���9��9/��93��9��9' �97�9V�9�9O �9���9��9���9���9���9\��9��9���9���9��9x   x   y��9F��9���9��9���9���9'��9���9���9q��9���9��9W��9A�9��9��9���9� �9��9���9�9^��9���9���9���9���9=��9���9��9���9x   x   ��9V��9���9;��9:��9��9L��9���9���97��9���9���9���9O��9m��9���9G��9W��9��9���9���9l��9&��9���9b��9���9��9:��9���9V��9x   x   P��9���9N��97��9^��9���9{��9���9��9��9���9��9��9���9���9��9:��9���9d��9d��9]��9���9��9��9���95��9���9���9��9!��9x   x   ���9P��9���9���9
��9L��9���9���9��9e��9���9T��9���9���9��9���9���9<��9���9R��9t��9<��9{��9���9��9��9���9���98��9���9x   x   9��98��9���9K��9P��9���9���9S��9r��9���9/��9���9��9���9v��9g��9��9]��9%��9_��97��9���9���9,��91��9b��9���9���9U��9���9x   x   5��9\��9
��9R��9���9���9d��9���9���9���9���9���91��9���9o��9r��9���9���9z��9���9V��9��9��9���9���9q��9 ��9x��9i��9���9x   x   ��9���9P��9���9���9h��9D��9z��9���9Z��9m��9���9<��9���9a��9g��9A��9���9!��9j��9;��9]��9��9S��9���9���9Q��9��9���9���9x   x   L��9|��9���9���9b��9A��9:��9n��9���9-��9���9���9���9X��9���93��9���9y��9���9���9���9w��9���9I��9y��9���9���9���9���98��9x   x   ���9���9���9U��9���9z��9v��9���9M��9<��9r��9���9~��9���9��9���9 ��9���9^��9{��9E��9���9l��9o��9(��9��9#��9���94��9S��9x   x   ���9��9��9q��9���9���9���9P��9���9���9���9j��9Q��9���9i��9���9���9#��9���9���96��9B��9���9���9��9���9p��93��9p��9
��9x   x   4��9��9f��9���9���9[��9(��9:��9���9{��9|��9���98��9���9?��9��9���9A��9���9���9���98��90��9���9���9w��9���9���9���9���9x   x   ���9���9���9+��9���9n��9���9s��9���9x��9-��9N��9)��9\��9x��9k��9v��9O��9���9@��9C��9���9���9z��91��9���9���9���9���9\��9x   x   ���9���9R��9���9���9���9���9���9l��9���9O��9���9���9+��9��9S��9���9���9h��9<��9��9���9R��9���9U��93��9���9(��9���9���9x   x   ���9��9���9��92��9B��9���9|��9R��98��9)��9���9���9��9���9O��9��9���9���9J��9}��9_��9G��9���9���9n��9���9���9���9���9x   x   O��9���9���9���9���9���9Z��9���9���9���9\��9+��9��9��9j��9q��9 ��9���9���9K��9���9���9x��9���9B��9P��9
��9B��9���9��9x   x   o��9���9	��9t��9k��9^��9���9��9g��9B��9x��9��9{��9i��9���9#��9���9!��9n��9���9\��9���9���98��9���9��9��9���9���9���9x   x   ���9��9���9n��9t��9j��94��9���9���9��9l��9Z��9Q��9r��9%��9^��9$��9���9��9���9���9���9���9���9v��9���9[��9D��9���9���9x   x   K��96��9���9��9���9>��9���9#��9���9���9q��9���9 ��9 ��9���9&��9���9���9��9'��9���9��9\��9���9���9���9��9��9s��9��9x   x   `��9���99��9]��9���9���9��9���9 ��9A��9Q��9���9���9���9"��9���9���9���9���93��9[��9���9���9���9���9\��9>��9r��9L��9��9x   x   ��9b��9���9#��9y��9 ��9���9^��9���9���9���9i��9���9���9j��9��9��9���9���9���9���9���9���94��9���9��9^��9���9���9`��9x   x   ���9g��9S��9c��9���9f��9���9z��9���9���9F��9A��9I��9K��9���9���9#��96��9���9���9���9\��9���9���9_��9���9���9?��9���9n��9x   x   ���9\��9v��9;��9S��98��9���9G��99��9���9B��9��9|��9���9]��9���9���9_��9���9���9@��9���9:��9��9���9���9-��9���9���9(��9x   x   f��9���9>��9���9��9\��9}��9���9?��96��9���9���9a��9���9���9���9��9���9���9\��9���9��9���9���9���9���9���9���9��9��9x   x   %��9��9z��9���9��9��9���9n��9���98��9���9O��9H��9x��9���9���9X��9���9���9���9;��9���9_��9|��9���9m��9���9���9���9}��9x   x   ���9%��9���9*��9���9P��9N��9n��9���9���9{��9���9���9���96��9���9���9���95��9���9��9���9x��9���9���9B��9���9���9p��9��9x   x   _��9��9��92��9���9���9x��9)��9��9���93��9S��9���9F��9���9u��9���9���9���9Y��9���9���9���9���9��9z��9c��9���9��9#��9x   x   ���93��9��9`��9r��9���9���9��9���9x��9���90��9t��9P��9��9���9���9Z��9��9���9���9���9n��9G��9z��9���9��9���9���9��9x   x   ��9���9���9���9��9V��9���9%��9r��9���9���9���9���9��9��9W��9��9=��9_��9���9,��9~��9���9���9b��9��9��9x��9���9���9x   x   6��9���9���9���9x��9��9���9���93��9���9���9'��9���9D��9���9D��9��9r��9���9?��9���9���9���9���9���9���9w��9H��9���9���9x   x   ���9��99��9V��9g��9���9���91��9n��9���9���9���9���9���9���9���9r��9F��9���9���9���9��9���9q��9��9���9���9���9���9'��9x   x   U��9%��9���9���9���9���95��9U��9	��9���9[��9���9���9��9���9���9��9��9a��9m��9&��9���9z��9��9&��9��9���9���9"��9:��9x   x   U��9���9��9���9��9��9Ð�9}��9���9���9��9���9ސ�9ɕ�9M��9��9j��9+��9���9T��9#��9���9Ւ�95��9���9��9���90��9�9ӏ�9x   x   ���9���9 ��9���9���9��9��9J��9c��9���9˗�9���9��9B��9ב�9��9ܒ�9��9�99��9:��9���9���9ސ�9Ɛ�9y��9@��9��9��9ِ�9x   x   ��9!��9;��9���9B��9���9���9���9ߑ�9���9ڕ�9���9���9ܒ�9ɗ�9��9���9̕�9ە�9i��97��94��9B��9_��9���9���9Ǌ�9ُ�9���9r��9x   x   ���9���9���9/��9���9��9��9u��9u��9ܖ�9��9��9O��9.��9���95��9���9d��9���9���9ϒ�9���9Ȓ�9���9W��9���9���9��93��9���9x   x   ��9���9A��9���9B��9<��9��9܏�9L��95��9���97��9���9Ւ�9���9Q��9~��9Δ�9��9��9g��9D��9���9|��9���9���9R��9ߎ�9���9 ��9x   x   
��9��9���9��9;��9���9���9���9��9f��9���9���9��9(��92��9���9���9ē�9��97��9���9"��9;��9���9$��93��9��9Y��9���9���9x   x   Ð�9��9���9��9��9���9��9q��9���9
��9t��90��9��9ϒ�9)��9���9{��9���9���9a��9��9���9���9t��9��9��9I��9=��9r��9g��9x   x   y��9H��9���9r��9��9���9q��9#��9���9��9$��9���9	��9)��9đ�9
��9��9��9,��9D��9ɑ�9ے�9��9���9���9:��9ҏ�9Ԑ�9$��9Q��9x   x   ���9`��9ܑ�9r��9N��9��9���9���9ڑ�9V��9��95��9֖�9œ�9J��9<��9̓�9͓�9���9{��9��9���9h��9t��9G��9���9���9-��9���9Ð�9x   x   ���9���9���9ݖ�98��9h��9��9��9X��9���9y��9��9u��9���9��9���9���9[��9��9?��9~��9���9U��90��9o��9��9}��9���9ɒ�9׌�9x   x   ��9ɗ�9ߕ�9��9���9���9u��9"��9��9u��9.��9]��9ԕ�9���9���9_��9[��9|��9;��9��9��9���9���92��9I��9)��9/��9���9���9��9x   x   ���9���9���9��98��9���9/��9���98��9 ��9[��9ۓ�9���9��9N��9���9���9ٕ�9|��9ϕ�9S��9��9���9l��9c��9ۓ�9��9��9��9��9x   x   ���9��9���9L��9���9��9��9��9ٖ�9w��9ו�9���9t��9]��9j��9g��9��9��9Ȑ�9���9ޕ�9���9|��9��9��9��9��9/��9ٖ�9I��9x   x   ȕ�9F��9��9-��9ؒ�9&��9ϒ�9(��9Ɠ�9���9���9��9`��9���9��9���9��9��9���9ƕ�9"��9��9���9���9D��9x��9۔�9���9��9^��9x   x   J��9֑�9ʗ�9���9���92��9)��9Ǒ�9J��9��9���9O��9k��9��9��97��9c��9��9Օ�9o��9@��9���9ו�9���9$��9���9��9��9���9�9x   x   ���9��9!��9.��9P��9���9���9��9:��9���9]��9���9c��9���95��9���9���9_��9���9ĕ�9e��9���9���9Ϙ�9��9*��9��9ԗ�9���9Ǖ�9x   x   e��9ޒ�9���9���9��9 ��9x��9��9Γ�9���9Z��9���9��9��9a��9���9���9Õ�9ٕ�9+��9ٖ�9���9.��9ɓ�9���9ܖ�9���9W��9	��9��9x   x   +��9��9ϕ�9b��9є�9œ�9���9��9ғ�9^��9w��9ܕ�9��9��9 ��9]��9���9���97��94��9���9��9���9���9��9 ��9���9��9<��9d��9x   x   ���9ɏ�9���9���9��9��9���9+��9���9��9<��9~��9Ő�9���9ו�9Ɨ�9ڕ�99��9!��9ї�9ח�9C��9v��9T��9ٕ�9��9�9��9���9l��9x   x   O��92��9h��9���9��9:��9c��9A��9|��9;��9
��9˕�9���9ƕ�9m��9ĕ�9-��96��9З�9ڏ�9���9ۘ�9���9���9��9Δ�9���9���9̔�9���9x   x    ��9;��94��9ɒ�9k��9��9��9Ƒ�9��9~��9��9W��9���9%��9@��9f��9ז�9��9ӗ�9���9���9���9ǖ�9ј�9���9ՙ�9���9ʓ�9j��9Ö�9x   x   ���9���93��9���9@��9 ��9���9ؒ�9���9���9���9��9���9��9��9���9���9��9D��9��9���9���9���9���9k��9w��9Ǔ�9B��9��9���9x   x   Ғ�9���9@��9ʒ�9���9>��9���9��9k��9U��9���9���9|��9���9ו�9���9-��9���9q��9���9Ȗ�9��9��9a��9���9
��9J��9���9B��9��9x   x   5��9ݐ�9\��9���9|��9���9o��9���9n��92��94��9n��9��9���9���9Ҙ�9Ǔ�9���9S��9���9՘�9��9b��9͓�9��9���9@��9 ��9r��9���9x   x   ���9ǐ�9���9T��9���9)��9��9���9K��9n��9I��9`��9��9@��9"��9���9���9��9ڕ�9��9���9j��9���9��9���9��9���9��9���9��9x   x   ��9z��9���9���9���95��9��9=��9���9��9-��9ٓ�9��9v��9���9.��9ݖ�9 ��9��9͔�9י�9v��9��9���9��9M��9��9j��9C��9��9x   x   ���9@��9Ǌ�9ߎ�9O��9��9H��9ҏ�9��9z��91��9��9��9ߔ�9��9��9���9 ��9���9���9���9Ǔ�9L��9=��9���9��9Q��9���9׍�9.��9x   x   .��9��9׏�9ߒ�9ގ�9U��99��9Ր�9*��9���9���9 ��92��9���9��9ԗ�9U��9��9��9~��9ʓ�9B��9���9!��9���9h��9Ð�9J��9/��9)��9x   x   �9��9���97��9���9���9p��9&��9���9͒�9���9��9ܖ�9��9���9���9
��9>��9���9̔�9j��9 ��9E��9u��9���9@��9׍�91��9��9���9x   x   Ϗ�9Ӑ�9n��9���9 ��9���9i��9S��9���9ӌ�9 ��9��9L��9_��9�9Õ�9��9h��9o��9���9���9���9��9ߑ�9��9��9+��9*��9���9���9x   x   lY�9\�9�\�9m]�9^�9�^�9�^�9 `�9�_�9]�9�^�9v_�9 d�96a�9�_�9pd�9�_�9�`�9d�9_�9^^�96]�9�_�9D`�9�^�9�^�97^�9,^�9�Z�9�[�9x   x   \�9�^�9�Z�9�]�9�_�9�_�9F`�9�]�9�^�9�Z�9�^�9�b�9Pb�9�^�9�c�9c�9i_�9bb�9�b�9X^�9n[�9_�9�\�9�`�9�_�9�_�9]�9�[�9�_�9�[�9x   x   �\�9�Z�9f[�9`a�9vZ�9[�9�\�9`�9�a�9�_�9�`�9�`�9O`�9c�9�d�9�b�9�_�9�`�9Ra�9�_�9�`�9`�9�\�9�Z�9�Z�9b�9�Z�9�Y�9)\�9�[�9x   x   i]�9�]�9`a�9a�9`�9l_�9�^�9{]�9Sa�9�[�9-^�9*^�9o^�98a�9�a�9o^�9�^�9�]�9�[�9"b�9�]�9�^�9�_�9�`�9�_�9�a�9S^�9�]�9P`�9�_�9x   x   ^�9�_�9zZ�9`�9zb�9I_�9n]�9!a�9�a�9N\�98e�9`�9�^�9�b�9^�9�_�9e�9�\�9a�9Fa�9?]�9'_�9"b�9�`�9�Z�9_�9�]�9�Z�9�W�9�[�9x   x   �^�9�_�9[�9p_�9I_�9�\�9r^�9�c�9�a�9f]�9�c�9�]�9ra�9~a�9^�9zc�9�]�9Nb�9�c�90^�9]�9�_�9�^�9�Z�9�_�9]_�9�\�9+Z�9�Y�9\�9x   x   �^�9D`�9�\�9�^�9n]�9o^�9`�9tc�9M_�9_�9d�9�`�9 b�9�`�9�c�9a_�9K^�9�c�9`�9�^�9i\�9�^�9]�9�_�9�^�9[�9ia�9�a�9�a�9r\�9x   x   "`�9�]�9`�9{]�9 a�9�c�9xc�9ub�9�c�9c�9�d�9da�9ka�9�d�9c�9d�9�b�96c�9�c�9^a�9/^�9�_�9�]�9=`�9�Y�9^�9l\�9	]�9V]�9>Y�9x   x   �_�9�^�9�a�9Ta�9�a�9�a�9L_�9zc�9ga�9�^�9Qa�9#^�9la�9�^�9�`�9�c�9_�98b�9aa�9?a�9Oa�9t^�9�_�9]b�9�\�9�a�9H]�9fa�9H]�9�b�9x   x   ]�9�Z�9�_�9�[�9N\�9f]�9_�9c�9�^�9�^�9{_�9u_�9~^�9)_�9:c�9_�9Y]�9Y\�9u\�95_�9�[�9:]�9�b�9�b�98a�9�b�9�b�90b�9�a�93b�9x   x   �^�9�^�9�`�9)^�96e�9�c�9d�9�d�9Qa�9|_�9�b�9{_�9�`�9�d�9�c�9
d�9e�9�]�9�`�9�^�9�]�9�]�9�[�9<^�9z_�9�_�9_�94]�9�\�9l^�9x   x   u_�9�b�9�`�9,^�9`�9�]�9�`�9ja�9&^�9w_�9z_�9�^�9Oa�9�`�9�]�9�_�9_�9a�9Nb�9*_�9�_�9lc�9ca�9a�9a�9`a�9�a�9�b�9lb�9�]�9x   x   �c�9Mb�9M`�9j^�9�^�9ka�9$b�9oa�9ha�9~^�9�`�9Na�9/b�9la�9�^�9�]�9�_�9�b�9Td�9`�9e_�9Qe�9jd�9De�9Dc�9�d�9�c�95d�9�a�9�`�9x   x   6a�9�^�9c�95a�9�b�9ua�9�`�9�d�9�^�9)_�9�d�9�`�9ma�9b�9�a�9�c�9�^�9�`�9�d�9;c�96a�9 _�9�`�95a�9�a�9Ja�92`�9�`�9�a�9Hd�9x   x   �_�9�c�9�d�9�a�9^�9^�9�c�9c�9�`�9:c�9�c�9�]�9�^�9�a�9�c�9�c�9�_�9�_�9`�9�d�9@d�9	b�9�f�9�g�9Cf�9�`�9�d�9�d�9�a�9`�9x   x   ud�9�c�9�b�9h^�9�_�9zc�9c_�9d�9�c�9_�9d�9�_�9�]�9�c�9�c�9d�9`�9Ld�9b�9{b�9_�9�`�9da�9Va�9b�9�^�9�b�9ub�9�b�9�_�9x   x   �_�9h_�9�_�9�^�9e�9�]�9L^�9�b�9_�9Y]�9e�9_�9�_�9�^�9�_�9`�9;b�9�c�9�b�9�e�9�f�9�e�9t_�9�d�9Nf�9�e�9b�9�c�9Nd�9�_�9x   x   �`�9`b�9�`�9�]�9�\�9Kb�9�c�92c�92b�9Y\�9�]�9a�9b�9�`�9�_�9Nd�9�c�9`�9,e�9�d�9g�9�b�9�c�9�f�9e�9Xe�9o`�9xc�9�b�9�_�9x   x   d�9�b�9Oa�9�[�9a�9�c�9`�9�c�9`a�9x\�9�`�9Pb�9Yd�9�d�9`�9b�9b�9*e�9�a�9�b�9Cf�9a�9�e�9*c�9	a�9 e�9Zb�9"b�9�a�9�d�9x   x   	_�9Y^�9�_�9"b�9Ia�9*^�9�^�9ca�9<a�99_�9�^�9,_�9`�9>c�9�d�9zb�9�e�9�d�9�b�9hk�9$g�9g�9�k�9�b�9�e�90e�9�b�9rd�9a�9�`�9x   x   e^�9q[�9�`�9�]�9@]�9
]�9h\�92^�9Na�9�[�9�]�9�_�9__�96a�9?d�9_�9�f�9 g�9Hf�9$g�9Nc�9g�9�e�9�f�9f�9N_�9�c�9b�9�`�9�^�9x   x   3]�9_�9�`�9�^�9%_�9�_�9�^�9�_�9m^�96]�9�]�9lc�9Me�9 _�9b�9�`�9�e�9�b�9a�9g�9g�9Za�9,c�9Te�9ea�9�a�9?_�9�d�9�a�9�]�9x   x   �_�9�\�9�\�9�_�9%b�9�^�9]�9�]�9�_�9�b�9�[�9ka�9id�9�`�9�f�9\a�9s_�9�c�9�e�9�k�9�e�9*c�9V_�9da�9f�9Da�9 d�98b�9�]�9�a�9x   x   I`�9�`�9�Z�9�`�9�`�9�Z�9�_�9>`�9ab�9�b�9;^�9a�9@e�99a�9�g�9Va�9�d�9�f�9-c�9�b�9�f�9Se�9ia�9h�9�a�9�d�9�a�9�\�9�a�9�c�9x   x   �^�9�_�9�Z�9�_�9�Z�9�_�9�^�9�Y�9�\�99a�9x_�9a�9Dc�9�a�9Cf�9b�9Rf�9e�9
a�9�e�9f�9ea�9f�9�a�92c�9�a�9�_�9b�9]�9�X�9x   x   �^�9�_�9b�9�a�9_�9^_�9~[�9 ^�9�a�9�b�9�_�9ca�9�d�9La�9�`�9�^�9�e�9We�9!e�90e�9L_�9�a�9Ea�9�d�9�a�9z^�9$c�9`a�9�]�9�\�9x   x   6^�9]�9�Z�9X^�9�]�9�\�9ja�9l\�9M]�9�b�9_�9�a�9�c�93`�9�d�9�b�9b�9n`�9Yb�9�b�9�c�9@_�9"d�9�a�9�_�9!c�9�\�9I]�9a�9�\�9x   x   .^�9�[�9�Y�9�]�9�Z�92Z�9�a�9]�9la�92b�92]�9�b�92d�9�`�9�d�9tb�9�c�9yc�9#b�9vd�9b�9�d�94b�9�\�9b�9`a�9I]�9�a�93Z�9�Z�9x   x   �Z�9�_�9)\�9M`�9�W�9�Y�9�a�9V]�9L]�9�a�9�\�9kb�9�a�9�a�9�a�9�b�9Od�9�b�9�a�9a�9�`�9�a�9�]�9�a�9!]�9�]�9a�92Z�9�W�9�_�9x   x   �[�9�[�9�[�9�_�9�[�9\�9t\�9;Y�9�b�90b�9m^�9�]�9�`�9Ed�9`�9�_�9�_�9�_�9~d�9�`�9�^�9�]�9�a�9�c�9�X�9�\�9�\�9�Z�9�_�9r]�9x   x   I)�9�*�9�(�9P'�9�+�9�(�9�*�96+�9=)�9%0�9�1�9E1�9B/�9�/�9�2�9�,�9�1�9�.�9p/�9�/�92�9�0�9;*�9�,�9�)�9�'�9O+�9�'�9�'�9�*�9x   x   �*�9;,�9l-�9�*�9|+�9�)�9�,�9�0�9�.�9�1�9)-�9{/�9�-�9�2�9e.�9F.�9�3�9~-�9�/�97.�9z1�9W.�9^.�9�,�9�*�9,�9�)�9�-�9�,�9�)�9x   x   �(�9q-�9�.�95&�9�/�90�9t-�9�,�9�-�9�0�9�.�9i-�9�.�9�/�9�&�9j/�9G.�9U-�9�.�9y/�9.�9A.�9�.�9m/�9�.�9�&�9G.�9�,�9s)�9�,�9x   x   Q'�9�*�94&�9&�9.�9<*�9-�9�,�9�+�9�.�9�2�9�.�93�90/�9�/�9�2�9�/�9[2�9h/�9�-�9+�9	,�9�)�9/�9&&�9&&�9�+�9�&�9,�9A,�9x   x   �+�9}+�9�/�9.�9�&�9N-�9=1�9�.�9�.�971�9�/�9t/�9m1�9�.�9v1�9h/�9a/�92�9�,�9�.�9)3�90-�9&�9.�9�/�9p*�9,�9�/�9�-�9�/�9x   x   �(�9�)�90�9=*�9J-�9�0�9�,�9G)�9&-�9�-�9�-�9�/�9G.�9�-�9 0�9�-�9�-�9�-�95*�9�+�9�/�9�.�9�)�9�/�9+�9a(�9�-�9-�9a,�9-�9x   x   �*�9�,�9p-�9-�9>1�9�,�9�,�9d+�9�/�9�-�9�-�9�-�9�/�9�-�9�-�9�.�9�.�9�+�99,�9�-�91�9,�9/�9�+�9h*�9@0�9�*�9L+�9}+�90�9x   x   5+�9�0�9�,�9�,�9�.�9G)�9c+�9-�9�,�9e,�9�)�9M/�9!/�9�)�9�+�9�,�9�-�9�*�9�)�9�.�9 -�9,,�9J0�9�+�9s1�9�/�9y,�9�,�9/�961�9x   x   >)�9�.�9�-�9�+�9�.�9%-�9�/�9�,�9=/�9�/�9f-�9�1�9�,�9�0�9:/�9`,�9�/�9.�9=-�9�+�9 /�9�-�9�)�9g+�9+�9|,�9`/�9B,�9�+�9�+�9x   x   #0�9�1�9�0�9�.�991�9�-�9�-�9h,�9�/�9�0�9�/�9�0�9#0�9�/�9�,�9�-�9/-�921�9Y1�9�.�9�1�9�0�9�0�9�-�9�,�9�+�9�+�9�,�9�,�9l1�9x   x   �1�9,-�9�.�9�2�9�/�9�-�9�-�9�)�9c-�9�/�9�,�9�/�9.�9&)�9,.�9}.�90�9)1�9[.�9�.�9F1�9�3�9V-�9�0�9E2�9�+�92�9�0�9!-�94�9x   x   E1�9|/�9l-�9�.�9p/�9�/�9�-�9E/�9�1�9�0�9�/�9�1�9�.�9.�9/�9w.�9�0�9�-�9�/�9�/�90�95/�9_,�90�9�-�9..�9�/�94-�9E.�9T/�9x   x   B/�9�-�9�.�93�9j1�9M.�9�/�9/�9�,�9#0�9.�9�.�90�9�-�9,3�9�1�9�-�9�-�9/�9�-�9�-�9�/�9�,�9�,�9i0�9c,�9#,�9�/�9J/�9�,�9x   x   �/�9�2�9�/�96/�9�.�9.�9�-�9�)�9�0�9�/�9*)�9.�9�-�9	.�9"/�91�9�2�9�/�9/�9M1�9�0�9�2�9\-�9�/�9�/�9.�93�9�/�9�1�9"/�9x   x   �2�9b.�9�&�9�/�9q1�9�/�9�-�9�+�9:/�9�,�9,.�9/�9)3�9/�9A&�9�-�9�2�9�1�9\.�9�0�9&0�9:3�9�/�9N/�9�.�9{2�9f1�9�/�9�.�991�9x   x   �,�9C.�9k/�9�2�9f/�9�-�9�.�9�,�9],�9�-�9{.�9y.�9�1�91�9�-�9�-�9U2�9/�9�.�9�1�9�/�9�3�9&/�9�/�9}4�9�.�9�1�9/�9�.�9>2�9x   x   �1�9�3�9I.�9�/�9[/�9�-�9�.�9�-�9�/�9,-�90�9�0�9�-�9�2�9�2�9P2�9g1�9�1�93�9�0�9 0�9�4�9�2�9u4�9�0�9D0�9H3�9�0�9�1�93�9x   x   �.�9}-�9U-�9]2�92�9�-�9�+�9�*�9.�901�9(1�9�-�9�-�9�/�9�1�9/�9�1�9u0�9H0�9�,�9�+�9�4�95�9�*�9�-�9u0�9�0�9'2�9p-�9<2�9x   x   n/�9�/�9�.�9j/�9�,�99*�9;,�9�)�9=-�9[1�9Y.�9�/�9/�9/�9U.�9�.�9#3�9J0�9�7�92�9�/�9X3�9�0�9�1�97�9�/�9�2�9�/�9�.�9�/�9x   x   �/�95.�9y/�9�-�9�.�9�+�9�-�9�.�9�+�9�.�9�.�9�/�9�-�9N1�9�0�9�1�9�0�9�,�92�9W0�9�.�9�-�9�0�9�1�9.�9�1�9~0�91�9�/�9�-�9x   x   2�9v1�9.�9+�9*3�9�/�91�9!-�9 /�9�1�9E1�9 0�9�-�9�0�9*0�9�/�90�9�+�9�/�9�.�9�.�9�.�9�/�9U+�9�-�9�0�9�/�9[1�9�.�9�/�9x   x   �0�9W.�9?.�9,�94-�9�.�9,�9/,�9�-�9�0�9�3�99/�9�/�9�2�983�9�3�9�4�9�4�9[3�9�-�9�.�913�9�4�9c6�9�3�93�9�2�9�.�9�.�923�9x   x   ?*�9a.�9�.�9�)�9&�9�)�9/�9I0�9�)�9�0�9V-�9^,�9 -�9^-�9�/�9'/�9�2�95�9�0�9�0�9�/�9�4�91�9�/�9�.�91.�9�-�9\,�9{.�9�0�9x   x   �,�9�,�9n/�9/�9.�9�/�9�+�9�+�9h+�9�-�9�0�90�9�,�9�/�9M/�9�/�9v4�9�*�9�1�9�1�9T+�9d6�9�/�9]/�9�/�93+�9m0�9�/�9�,�9+�9x   x   �)�9�*�9�.�9)&�9�/�9+�9i*�9r1�9+�9�,�9G2�9�-�9l0�9�/�9�.�9|4�9�0�9�-�97�9.�9�-�9�3�9�.�9 0�9�0�9e.�9Q2�9+-�9,�90�9x   x   �'�9,�9�&�9%&�9t*�9e(�9C0�9�/�9z,�9�+�9�+�9/.�9b,�9�.�9}2�9�.�9E0�9w0�9�/�9�1�9�0�93�90.�96+�9d.�9�*�9,�9X+�9�/�91�9x   x   L+�9*�9E.�9�+�9,�9}-�9�*�9y,�9]/�9�+�92�9�/�9 ,�93�9i1�9�1�9K3�9�0�9�2�9}0�9�/�9�2�9�-�9l0�9O2�9,�9�/�9�,�9*�9$.�9x   x   �'�9�-�9,�9�&�9�/�9�,�9L+�9�,�9@,�9�,�9�0�98-�9�/�9�/�9�/�9/�9�0�9&2�9�/�91�9[1�9�.�9a,�9�/�9--�9W+�9�,�9,�9�,�9e/�9x   x   �'�9�,�9p)�9,�9�-�9^,�9+�9/�9�+�9�,�9-�9E.�9N/�9�1�9�.�9�.�9�1�9o-�9�.�9�/�9�.�9�.�9u.�9�,�9,�9�/�9*�9�,�9.�9,�9x   x   �*�9�)�9�,�9A,�9�/�9-�90�971�9�+�9q1�94�9U/�9�,�9$/�961�9>2�9"3�9;2�9�/�9�-�9�/�933�9�0�9+�9�0�9
1�9(.�9g/�9,�9�-�9x   x   �9���9��9-��9,��9���9���9J��9��9���9���9�9G��9���9d��9r��9!��9=��9���9��9���9��9
 �9���9���9���9��9���9���9���9x   x   ���9���9Y��9���9���9	��9Q��9���9q��9���9���9���9n��9%��9��9��9���9x��9���9���9���9���9���9��9���9���9��9s��9q��9b��9x   x   ��9R��9%��9��9T��9c��9,��9���9���9f��9���9' �9o��9���9�9$��9���9. �9��9���9��9���9���9���9���9���9���9\��9��9��9x   x   .��9���9~��9���9���9���9b��9�9���9���9���9���9���9���9L �9���9���96��9#��9���9���9M��9���9���9j��9���9���9Q��9#��9\��9x   x   .��9���9T��9���9���9���9���9���9��9Z��9���9���9���9c��9e��9h��9���9���9T��9���9��9j��9���9=��9���9���9���9
��9���9���9x   x   ���9��9g��9���9���9?��9C��9m��9���9���9���9� �9��9���9� �9��9i��9���9���9P��9���9���9���9���9���9Z��9���9T��9t��9���9x   x   ���9Q��9.��9g��9���9D��9��9���9��9$�9��9���9D��9  �9'��9A�9� �9%��9��9]��9���9��9���9���9���9K��9&��9���9��9D��9x   x   J��9���9���9�9���9n��9���9)��9���9l��9Y�9���91��9�9���9\��9���9��9���9���9� �9 ��9��9C��97��9���9��9���9<��9���9x   x   	��9o��9���9���9��9���9��9���9S��9
 �9���9S��9���9�9���96��9��9���9���9���9'��9{��9���9F��9� �9,��9���9V��9v �9T��9x   x   ���9���9f��9���9X��9���9!�9i��9 �9S��9���9;��9���9Z��9���9� �9��9��9� �9���9���9���9���9���9���9���9���9���9Q��9���9x   x   ���9���9���9���9���9���9��9_�9���9���9���9���9]��9� �9���9���9Z��9f��9#��9���9���9)��9j �9.��9���9>�9[��9���9���9��9x   x   � �9���9% �9���9���9� �9���9���9X��9:��9���9p��9��9� �9���9���9� �9} �9���9���9F��9��9��9���9W��9)��9���9� �9.��9��9x   x   H��9p��9m��9���9���9��9A��95��9���9���9[��9��9���9|��9���9���9��9���9���9��9o�9u��9c �9�9��9/�9� �9~��9� �9+��9x   x   ���9#��9���9���9^��9���9 �9�9�9X��9� �9� �9��9��9���9��9���9���99��9���9O��9 �9��9
�9�9E�9?��9N��9��9���9x   x   g��9��9�9H �9d��9� �9$��9���9���9���9���9���9���9���9��9?�9N��9B �9��9���9���9Z��9���9 �9#��9���9V��9%��9;�9Y��9x   x   r��9��9#��9���9j��9��9?�9\��98��9� �9���9���9���9��9A�9��9���99��9��9� �9�9��9��9��9���9��9� �9��9\�9���9x   x   #��9���9���9���9���9l��9� �9���9��9��9X��9� �9��9���9O��9���9���9���9Q��9'�9��9���9���9A��9��9 �9���9a��9���9���9x   x   =��9}��9/ �95��9���9���9#��9
��9���9��9f��9� �9���9���9H �99��9���9��9���9S�9��9g��9-��9�9��9[��9��9b��9���9� �9x   x   ���9���9��9��9Z��9���9��9���9���9� �9!��9���9���9;��9��9��9M��9���9Q �9J�9��9��9��9��91 �9���9*��9��9/�9Q��9x   x   ��9���9���9���9���9X��9a��9���9���9���9���9���9��9���9���9� �9"�9S�9H�9���9��95�9���9�9`�9��99��9��9I��9� �9x   x   ���9���9��9���9��9���9���9� �9'��9���9���9I��9p�9J��9���9�9��9��9��9��9b�9��9@�9�9���9��9_��9)��9'�9���9x   x   ��9���9���9Q��9g��9���9��9���9���9���9(��9��9u��9 �9Y��9��9���9n��9��99�9��9��9W��9���9C��9���9��9y��9���9H��9x   x    �9���9���9���9���9���9���9��9���9���9i �9��9h �9��9���9��9���90��9��9���9=�9U��9���9]�9���9��9m�9� �9 �9���9x   x   ���9��9���9���9B��9���9���9D��9A��9���92��9���9�9�9 �9��9=��9�9 �9"�9�9���9Z�9���9��9���9���9���9���9v��9x   x   ���9���9���9j��9���9���9���9=��9� �9���9���9T��9��9�9 ��9���9��9��92 �9d�9���9E��9���9��97 �9���9���9���9��9���9x   x   ���9���9���9���9���9V��9J��9���9-��9���9?�9%��91�9F�9���9��9 �9Z��9���9��9��9���9��9���9���9��9���9���9���9���9x   x   ��9��9���9���9���9���9'��9��9���9���9\��9���9� �9<��9Y��9� �9���9��9,��9;��9_��9!��9l�9���9���9���9� �9���9A��9I��9x   x   ���9q��9a��9O��9��9T��9���9���9W��9���9���9� �9���9N��9!��9��9`��9a��9��9��9-��9y��9� �9���9���9���9���9���9S��9y��9x   x   ���9s��9��9#��9���9r��9��9A��9w �9T��9���9)��9� �9��9=�9[�9���9���9,�9G��9'�9���9 �9���9��9���9A��9Q��9���9|��9x   x   ���9`��9��9[��9���9���9A��9���9Q��9���9��9 ��9$��9���9a��9���9���9� �9T��9� �9���9H��9���9x��9���9���9C��9t��9{��9(��9x   x   ���9H��9&��9I��9_��9���9��9Q��9���9���9O��9 ��9-��9f��9��9D��9���9J��9��9v��9���9���9���9���9;��9s��9���9���9u��91��9x   x   G��9���9���9���9���9���9 ��9U��9���9r��9���9���9���9���9���9���9���9���9���9���9>��9���9���9���9���9���9 ��9���9���9C��9x   x   )��9���9���9���9��9���9���9���9��9���9��9���9*��9��9!��9���9���9
��9���9���9+��9u��9F��9��9]��9@��9&��9��9���9���9x   x   K��9���9���9���9V��9���9/��9���9���9 ��9W��9v��9���91��9$��9b��9z��9���9���9W��9���9V��9U��9���97��9a��9T��9���9���9���9x   x   `��9���9��9X��9��9���9��9���9?��9���9���9���9��9���96��9Z��9_��9��9��9���9��9���9���9��9���9��9���9u��9���9-��9x   x   ���9���9���9���9���9���9��9���9���9���91��9	��9;��9��9���9���9T��9��9E��9��9U��9���9��9��9���9���9��9#��9j��9u��9x   x   ��9��9���90��9��9��9r��9B��9��9���9(��9T��9_��9���9���9���9��9M��9���9���9p��9)��9��9���91��9���9&��9?��9	��9���9x   x   Q��9V��9���9���9���9���9@��9���9���9���9^��9���9
��9���9'��9���9A��9���9���9��9 ��9���9���9I��9���9o��9o��9���9/��9i��9x   x   }��9���9��9���9?��9���9$��9���9���9���9 ��9}��9��9���9e��9��9Z��9���9���94��9l��9&��9@��9��9}��9���9���9���9���9e��9x   x   ���9o��9���9!��9���9���9���9���9���9 ��9a��9���9I��9U��9���94��9+��9h��9���9���9E��98��9q��9���9���9��9���94��9a��9���9x   x   Q��9���9��9X��9���9-��9(��9[��9��9c��9���9���9��9���9a��9|��9���9e��9p��9���9���9���9���9:��9���9���9e��9���9g��9���9x   x   ���9���9���9w��9���9
��9T��9���9t��9���9���9���9���9{��9���9���9���9Y��9���9���9���9���9���9���9��9q��9���9���9R��9���9x   x   +��9���9-��9���9��96��9`��9
��9��9Q��9��9���9���9���9��9��9���9���9���9-��9���9L��9���9���9���9 ��9U��9*��9Y��9P��9x   x   h��9���9}��95��9���9��9���9���9���9V��9���9}��9���9���9\��9S��9���9���9���9u��9���9���9P��9���9/��9C��9H��9���9���9��9x   x   ��9���9��9)��96��9���9���9*��9d��9���9a��9���9��9Z��9���9B��9���9 ��9���9���9���9���9���9d��9��9��9H��9���9(��9A��9x   x   ?��9���9���9e��9V��9���9���9���9!��96��9}��9���9��9T��9@��9i��9��9$��9���9���9���9;��96��9���9���9]��9���9y��9���9���9x   x   ���9���9���9}��9a��9R��9���9C��9T��9(��9���9���9���9���9���9	��9���9���9��9��9���9v��9d��9-��9}��9W��9��9���9���9"��9x   x   G��9��9	��9���9��9��9T��9���9���9f��9j��9[��9���9���9��9#��9���9��9���9���9���9_��9���9���9���9���9a��9J��9O��9r��9x   x   ��9���9���9���9��9B��9���9���9���9���9m��9���9���9���9���9���9��9���9��9y��9���9���9���9i��9���9���9K��9���9��9���9x   x   w��9���9���9X��9���9��9���9��97��9���9���9���9/��9t��9���9��9��9���9w��9S��9���9���9k��9���9���9��9���9���9%��9���9x   x   ���9<��9,��9���9��9P��9q��9���9h��9B��9���9���9���9���9���9���9���9��9���9���9���9���9P��9b��9���9���9��9F��9���9��9x   x   ���9~��9x��9Y��9���9���9.��9���9&��96��9���9���9Q��9���9���9<��9t��9b��9���9���9���9��9���9Y��9 ��9��9��9���9���9���9x   x   ���9���9F��9Q��9���9��9��9���9@��9t��9���9���9���9K��9���94��9`��9���9���9j��9L��9���94��9���9s��9��9���9��9}��9g��9x   x   ���9���9��9���9��9��9���9K��9��9���9<��9���9���9���9c��9���9/��9���9j��9���9c��9[��9���9���9���9��9���9���9��9���9x   x   ?��9���9`��93��9���9���93��9���9~��9���9���9��9���93��9��9���9~��9���9���9���9���9��9u��9���9���9|��9j��9���9��9���9x   x   r��9 ��9C��9a��9��9��9���9f��9���9��9���9t��9��9C��9��9Z��9Y��9���9���9��9���9���9��9��9���94��9g��9���9���9q��9x   x   ���9��9(��9V��9���9��9'��9n��9���9��9e��9���9V��9G��9F��9���9��9d��9J��9���9��9��9��9���9n��9d��9���9��9"��94��9x   x   ���9���9��9���9r��9!��9B��9���9���91��9���9���9+��9���9���9|��9���9L��9���9���9C��9���9��9���9���9���9��9���9R��9���9x   x   x��9���9���9���9���9n��9��9)��9���9b��9l��9R��9Y��9���9$��9���9���9R��9���9)��9���9���9}��9��9��9���9 ��9W��9���9��9x   x   2��9G��9���9���9/��9z��9���9g��9c��9���9���9���9P��9x��9<��9���9��9p��9���9���9!��9���9d��9���9���9s��96��9���9��9���9x   x   Ф�9���9˜�97��9���9���9���9��9��9K��9D��9���9��9d��9|��9���9;��9��9$��9.��9��9ŝ�9��9���9��9���9?��9���9��9���9x   x   ���9��9i��9L��9���9��9o��9j��9#��9��9X��9���9���9���9���9 ��9��9���9���9)��9��9��9Ο�9��9��9o��9���9l��9���9B��9x   x   ̜�9p��9V��9ڝ�9���9���9?��9��9��9H��9���9���9��9ť�9$��9���9��9��9+��9��9@��9���9\��99��9{��9)��9a��9��9���9A��9x   x   5��9O��9ם�9:��9��9��9~��9L��9���9��9s��9��9g��9۠�9���9O��9���9[��9��9*��9j��9��9ԟ�9���9H��9���9���9��9.��9���9x   x   ���9���9���9��95��9+��9��9K��9��9���9��9���9���9u��9��9���9<��9ء�9О�9W��9E��9���9��9-��9���9���9���9˟�9F��9r��9x   x   ���9��9���9��9)��9u��9*��9M��9���9n��98��9T��9y��98��9>��9���9}��9A��9��9T��99��9b��90��9���9e��9���9���9G��9��9	��9x   x   ���9q��9>��9���9��9)��9���9��9���9���9M��9#��9���9j��9f��9/��9��9���9���9}��91��9j��9���9���9ҟ�9"��9A��9��9ʟ�9���9x   x   ��9o��9��9N��9O��9M��9��9���9A��9���9���9���9J��9���9ˡ�9ܠ�9��9���9���9��9y��9Q��9��9Y��9>��9���9/��9��9���9+��9x   x   ��9(��9��9���9z��9���9z��9=��9¢�9��9-��9֡�9R��9Ѥ�9���9ٟ�9D��9��9��9���9���9n��9М�9���9V��9���9D��9|��9;��9���9x   x   K��9��9F��9��9���9q��9���9���9��9˦�9���9D��9���9��9 ��9&��9���9ʠ�9%��9s��9���9���9v��9���9۠�9@��9&��9~��9��9���9x   x   E��9X��9���9u��9��99��9M��9���92��9���9t��9ؠ�9��9��9h��9f��9���9@��9���9��9���9���9��9���9Q��9���9٢�9T��9B��9i��9x   x   ���9���9���9��9���9U��9$��9���9ء�9F��9ՠ�9���9/��9��9���9��9��9"��9���9֠�9A��9u��9Ǡ�9���9���9��9ԣ�9���9���9��9x   x   ��9���9��9a��9���9z��9���9M��9V��9���9��9/��98��9��9e��9���9"��9���9���9��9���9��9;��9���9ף�98��9ܡ�9ݡ�9��9Ρ�9x   x   b��9���9ĥ�9٠�9t��99��9j��9���9Ԥ�9��9��9��9��9���9	��9���9\��9��9ģ�9���9���9=��9Ϡ�9(��9���9?��9��9��9���9'��9x   x   |��9���9#��9���9��9A��9h��9ˡ�9���9��9i��9���9g��9��9��9ӟ�9%��9=��9���9���9j��9Σ�9t��9��9���9Ѣ�9c��9��9;��9��9x   x   ���9"��9���9M��9���9���92��9ڠ�9۟�9'��9f��9��9���9���9џ�9C��9��9ˡ�91��9���9���98��9{��9��9y��9V��95��9=��9\��9V��9x   x   ;��9	��9��9���9<��9���9��9 ��9J��9���9���9��9"��9^��9%��9��9q��9���9��9)��9��9���9���9���9���9#��9J��9��9 ��9i��9x   x    ��9���9��9[��9ء�9C��9���9���9��9ʠ�9A��9"��9���9��9<��9̡�9���9e��9q��9���9v��9��9i��9���9���9_��9	��9}��9:��9���9x   x   &��9���9-��9��9О�9��9���9���9
��9%��9���9���9���9ƣ�9���91��9��9n��9��9a��9���9���9��9ĥ�9��9���9;��9���9G��9��9x   x   .��9)��9��9(��9X��9T��9��9��9���9u��9��9Ҡ�9��9���9���9���9*��9���9d��9K��9���9��9A��9���9ʣ�9A��9���9,��9x��9*��9x   x   ��9��9?��9i��9H��9<��91��9v��9���9���9���9A��9���9���9g��9���9��9q��9���9���9���9ç�9E��9Ν�9���9��9R��92��9Ƞ�92��9x   x   Ɲ�9"��9���9��9ɞ�9j��9g��9U��9p��9���9���9u��9��9>��9ϣ�9:��9���9���9���9��9§�9���9e��9���9Ǥ�9���9���9D��92��9#��9x   x   ��9П�9Z��9П�9��9,��9��9��9Ϝ�9u��9��9Ơ�99��9Ҡ�9u��9~��9���9i��9��9@��9I��9l��9G��9���9��9w��9���9���9٠�9���9x   x   ���9��9:��9���91��9���9���9V��9 �9���9���9���9���9)��9��9��9���9���9ť�9���9̝�9���9~��9ߠ�9���9��9D��9Z��9^��9��9x   x   ��9��9w��9H��9���9a��9џ�9=��9X��9ޠ�9T��9���9֣�9���9���9x��9���9���9��9ˣ�9���9Ĥ�9��9���9[��9a��9ܣ�9,��9���9*��9x   x   ���9m��9(��9���9���9���9)��9���9���9?��9���9��93��9@��9Ӣ�9V��9#��9_��9���9@��9��9 ��9u��9	��9\��9&��9	��9w��9��9��9x   x   ?��9��9a��9���9���9���9D��9/��9C��9$��9آ�9գ�9١�9��9d��94��9D��9��9:��9���9U��9���9���9B��9٣�9��9ƣ�9a��9j��9ȟ�9x   x   �9q��9��9��9ϟ�9E��9��9��9���9���9T��9���9ޡ�9��9��9;��9��9z��9���9*��9.��9F��9���9[��9-��9y��9d��9k��99��9;��9x   x   ��9���9���92��9H��9��9͟�9���9:��9��9@��9���9��9���9=��9_��9 ��9<��9K��9y��9Ơ�94��9ܠ�9_��9���9��9j��97��9��9��9x   x   ���9A��9C��9���9q��9��9��9,��9���9���9g��9��9ϡ�9)��9��9V��9f��9���9��9*��90��9 ��9���9!��9,��9��9Ɵ�96��9��9���9x   x   l�9�o�9Tv�9�u�9ls�9�u�9�t�9/r�9�u�9�u�9�s�9u�9�u�9bs�9bv�9Pt�9�u�9t�9yv�9�u�9,s�9�t�9�u�9|r�9�t�9u�9t�9v�9�u�9�o�9x   x   �o�9[n�95q�9�o�9�r�9�r�9�q�9�w�9�u�9hu�9Mt�91x�9�x�9�s�9 w�9:x�9�s�9�w�9�w�9�s�9fv�9�v�9�v�9Cq�9qs�9�r�9Go�9+q�9�n�9-p�9x   x   Pv�91q�9�p�9s�9�u�93p�9�p�9�q�9't�9ut�9+p�9�v�9s�9t�9z�9s�9�s�9Aw�9�p�9�t�9�r�9q�9)r�9p�9�u�9Ss�9q�9Jq�9Ku�9Nw�9x   x   �u�9�o�9s�9Mr�9s�9v�9�u�9}s�9ax�96t�9�u�9[x�9�q�9u�9u�9~r�9x�9�t�9�s�9�x�9�t�9�u�9^u�9�r�9Er�9s�9Co�95v�9Ru�9=t�9x   x   fs�9�r�9�u�9s�9�w�9�v�9�t�9Su�9s�9Us�9�t�9�w�9{v�9ft�9�v�9vv�9�u�9�s�9�r�9Gu�9/t�9-v�9�x�9�s�9Fu�9Us�9^s�9�s�94n�9�t�9x   x   �u�9�r�96p�9v�9�v�9^i�9ss�9Ws�9�r�9�u�9}r�9Fv�9�s�9?s�9�v�9s�9�t�9�r�9}s�9s�9�j�9]v�9�t�9cp�9�r�9Pu�9ut�9�v�9+v�9�s�9x   x   �t�9�q�9�p�9�u�9�t�9rs�9?y�9�p�9�t�9�u�9v�9�u�9�t�9�u�9�u�9`u�9�u�9Gp�9�y�9?s�9�s�9�v�9�q�9�q�9�t�9�r�9�p�9�{�9�p�9js�9x   x   0r�9�w�9}q�9�s�9Pu�9\s�9�p�9`r�9�s�9(r�9�s�9t�9�t�9�s�9yr�9t�9�q�9�p�9Cs�9�u�9�s�9�p�9�v�9�q�9�t�9�q�9u�9~u�9�q�9�s�9x   x   �u�9�u�9't�9^x�9s�9�r�9�t�9�s�9t�9yt�90s�9:v�9�r�9�t�9Ms�9Vs�9'v�9/r�9s�9�x�9_s�9>v�9�v�9�s�9�s�9v�9w�9=u�9t�9�t�9x   x   �u�9ku�9wt�98t�9Ws�9�u�9�u�9"r�9wt�9�o�9�t�9�t�96p�9�t�9s�9$u�9�t�9*t�9ls�9�t�9v�9rt�9`x�9Gw�9�r�9�s�9At�9Ss�9�v�9x�9x   x   �s�9Lt�9&p�9�u�9�t�9}r�9v�9�s�9,s�9�t�9�x�9�t�9�r�9�s�9�u�9>s�9(u�9}u�9�p�9�s�9�s�9Lr�9u�9�s�9u�9�x�9Ut�97s�9�u�9]r�9x   x   u�92x�9�v�9\x�9�w�9Gv�9�u�9t�96v�9�t�9�t�97v�9�t�9Bv�9�v�9w�9�w�9w�9�w�9�t�9�t�9�v�9�t�9p�9Vs�9�s�9q�9Au�9yv�9�s�9x   x   �u�9�x�9s�9�q�9|v�9�s�9�t�9�t�9�r�90p�9�r�9�t�9St�9�s�9�u�9!s�9�s�9x�9w�9Tu�9Iu�9�u�9�v�9t�9�t�9
s�9�u�9�t�9�v�9�v�9x   x   es�9�s�9t�9u�9et�9As�9�u�9�s�9�t�9�t�9�s�9?v�9�s�9�t�9�t�9�r�9�s�9s�9�r�9�w�9�r�9Pv�9�u�9�s�9�t�9�v�9-w�9�r�9�u�9%s�9x   x   fv�9�v�9z�9
u�9�v�9�v�9�u�9tr�9Ps�9s�9�u�9�v�9�u�9�t�9�z�9�w�9�v�9{v�9u�91v�9�u�9�u�9Jr�9x�9/q�9�t�9>u�9w�9�u�9�v�9x   x   Pt�9:x�9s�9�r�9{v�9s�9_u�9t�9Vs�9!u�9>s�9w�9s�9�r�9�w�9�r�9�v�9v�9�t�90u�9�t�9�q�9�z�9�z�9�r�9�u�9�t�9�t�9\u�9	v�9x   x   �u�9�s�9�s�9x�9�u�9�t�9�u�9�q�9(v�9�t�9(u�9�w�9�s�9�s�9�v�9�v�94t�9�v�9w�9w�90x�9�v�9s�9w�9�v�9�w�9�v�9�v�9�u�9v�9x   x   t�9�w�9Bw�9�t�9�s�9�r�9Ip�9~p�9-r�9(t�9{u�9w�9
x�9s�9v�9~v�9�v�9�w�9�r�9t�9�y�9u�9?t�9�y�9�t�9�r�9'x�91v�9�u�9w�9x   x   xv�9�w�9�p�9�s�9�r�9~s�9�y�9>s�9
s�9ns�9�p�9�w�9�v�9�r�9u�9�t�9w�9�r�9ts�9�w�9ft�9�x�9�t�9jx�9�r�9xr�9<w�9�t�9�u�9Xr�9x   x   �u�9�s�9�t�9�x�9Du�9	s�9As�9�u�9�x�9�t�9�s�9�t�9Pu�9�w�91v�93u�9w�9t�9�w�9pq�9�r�9js�9p�9gw�9�u�9yv�9Ou�9kv�9w�9�u�9x   x   )s�9jv�9�r�9�t�9/t�9�j�9�s�9�s�9as�9v�9�s�9�t�9Ju�9�r�9�u�9u�93x�9�y�9et�9�r�9�q�9�r�9�u�9y�9Aw�9�u�9Fu�9�r�9sv�9jt�9x   x   �t�9�v�9q�9�u�9$v�9Yv�9�v�9�p�9<v�9st�9Lr�9�v�9�u�9Nv�9~u�9�q�9�v�9u�9�x�9js�9�r�9 x�9@t�9!w�9�r�9�t�9w�9[u�9�u�9�r�9x   x   �u�9�v�90r�9`u�9�x�9�t�9�q�9�v�9�v�9^x�9u�9�t�9�v�9�u�9Jr�9�z�9s�9@t�9�t�9p�9�u�9@t�9�s�9Iz�9�q�9v�9"v�9�t�9v�9�w�9x   x   �r�9Cq�9p�9�r�9�s�9dp�9�q�9r�9�s�9Kw�9�s�9p�9t�9�s�9x�9�z�9	w�9�y�9hx�9ew�9y�9#w�9Kz�9�x�95t�9�s�9�p�9ys�9;v�9�t�9x   x   �t�9ns�9�u�9Dr�9Cu�9�r�9�t�9�t�9{s�9�r�9u�9Ts�9�t�9�t�90q�9�r�9�v�9�t�9�r�9�u�9Cw�9�r�9�q�99t�9Ct�9�s�9Qt�9cs�9�s�9�s�9x   x   u�9�r�9Xs�9s�9Xs�9Qu�9�r�9�q�9
v�9�s�9�x�9�s�9s�9�v�9�t�9�u�9�w�9�r�9ur�9uv�9�u�9�t�9v�9�s�9�s�9�x�99t�9�u�9�q�9�s�9x   x   t�9Fo�9q�9Co�9bs�9st�9�p�9u�9w�9Ft�9St�9q�9�u�9+w�9Au�9�t�9�v�9)x�9Dw�9Nu�9Eu�9w�9v�9�p�9St�9:t�9bv�9�u�9�p�9�s�9x   x   v�9)q�9Kq�91v�9�s�9�v�9�{�9�u�9:u�9Ss�98s�9Au�9�t�9�r�9w�9�t�9�v�91v�9�t�9iv�9�r�9`u�9�t�9xs�9bs�9�u�9�u�9�z�9�v�9�s�9x   x   �u�9�n�9Nu�9Ju�94n�9-v�9�p�9�q�9t�9�v�9�u�9{v�9�v�9�u�9�u�9Zu�9�u�9�u�9�u�9w�9pv�9�u�9 v�9:v�9�s�9�q�9�p�9�v�9�n�9�t�9x   x   �o�9-p�9Mw�97t�9�t�9�s�9gs�9�s�9�t�9x�9^r�9�s�9~v�9#s�9�v�9v�9v�9w�9Wr�9�u�9ht�9�r�9�w�9�t�9�s�9�s�9�s�9�s�9�t�9�w�9x   x   O�9�J�9rH�9\J�9�D�9�I�9I�9�G�9�H�9rJ�9NL�9G�9�J�99L�9�H�9�I�9rH�9�M�9oJ�9/H�9nK�9�I�9�H�9�F�9�I�9FJ�9cE�9~J�9�G�9�J�9x   x   �J�9{J�9�J�9I�9G�9�H�9!M�9(H�9�E�9�G�9�M�9�D�9�I�9/J�9G�9NH�9�H�9�H�9E�9�L�9I�9�E�9?I�9	M�9H�9�F�9�H�9vJ�9�J�9L�9x   x   uH�9�J�9I�9L�9-G�9�K�9�J�9QJ�9�I�9�H�9L�9eF�9�I�9�H�9�H�9�H�95K�9G�9fK�9ZI�9I�9I�9�J�93L�9�G�9L�9{I�9�J�9�F�9�B�9x   x   bJ�9I�9
L�9�H�9cH�9�F�95G�9cI�9�H�91I�9@H�9�J�99H�9�I�9�H�9_H�9�I�9�G�9J�9jG�9OK�9�G�9�F�9H�9_H�9QL�9�G�9�K�9�H�9jG�9x   x   �D�9G�9.G�9dH�9F�9�G�9�K�9DG�9�K�9�J�9BI�9�K�9�G�92M�9I�9+K�9iJ�9�J�9L�9G�9�I�9�G�9aF�9�H�9�F�9�G�9�D�9RG�9 H�9QH�9x   x   �I�9�H�9�K�9�F�9�G�9�M�9_K�9G�9�K�9nJ�9vJ�9F�9�I�9qI�9�E�9�J�9�I�9,K�9PH�9�K�9O�93G�9QF�9OL�9�G�9aJ�9I�9PF�9<F�9�H�9x   x   I�9 M�9�J�92G�9�K�9`K�9�H�9iJ�9�G�9UG�9�G�9&H�9L�9�G�9&H�9{F�9�I�9J�9H�9�J�9�J�9fH�9J�9�M�9�H�9K�9=I�9EG�9�H�9�K�9x   x   �G�9(H�9VJ�9aI�9DG�9{G�9gJ�9O�9L�9�I�9^L�9dG�9^H�9=L�9�I�9�K�9�M�9K�9*H�9�G�9^I�9`J�9(H�9�G�9�E�9\K�9E�9�E�9~K�90E�9x   x   �H�9�E�9�I�9�H�9�K�9�K�9�G�9L�9K�9'J�9�N�9�H�9�M�9�I�9�K�9L�9�H�9K�9SK�9I�9mH�9PF�9�H�9G�9�J�9�K�9B�9LK�9�J�9^G�9x   x   rJ�9�G�9�H�9/I�9�J�9jJ�9VG�9�I�9(J�9�H�9�I�9zI�9J�9�I�9�I�9vG�9�I�9�K�96H�9�I�9�H�9�I�9,I�9�G�9MI�9�G�9�G�9�I�9H�9H�9x   x   RL�9�M�9L�9BH�9BI�9sJ�9�G�9cL�9�N�9�I�9�I�9�I�9�M�9�L�9�G�9�J�9UI�9�H�9�K�9>L�9,L�9�I�9�F�9	J�9BI�9�K�9;I�9�H�9�G�9	J�9x   x   	G�9�D�9iF�9�J�9�K�9F�9(H�9fG�9�H�9}I�9�I�9�H�9lH�99H�96F�9�L�9�H�9~F�9�E�9H�9J�9OJ�9�J�9L�9�I�9�I�9�L�9�J�93J�9�I�9x   x   �J�9�I�9�I�96H�9�G�9�I�9L�9^H�9�M�9J�9�M�9mH�9�J�9:J�9�F�9�I�9jK�9�H�9]J�9H�9�H�9�H�9�H�9M�9~J�9�K�9-I�9_H�9,I�9�I�9x   x   8L�90J�9�H�9�I�91M�9sI�9�G�9?L�9�I�9�I�9}L�9<H�9;J�9HN�9"I�9 G�9�I�9�L�9�I�9�H�9K�9MG�9lJ�9�I�91K�9�J�9LG�9�K�9LG�9�H�9x   x   �H�9G�9�H�9�H�9I�9�E�9-H�9�I�9�K�9�I�9�G�95F�9�F�9$I�9�I�9�G�9�H�9&I�9�G�9M�9PL�9M�9RJ�9�G�9oI�9�L�9�K�9�M�9GI�9�I�9x   x   �I�9KH�9�H�9\H�9*K�9�J�9~F�9�K�9 L�9wG�9�J�9�L�9�I�9�F�9�G�9I�9�J�9�I�9{I�9&H�9L�9mI�9 L�9�K�9J�9�L�99G�9�H�9�H�9�J�9x   x   sH�9�H�98K�9�I�9nJ�9�I�9�I�9�M�9�H�9�I�9YI�9�H�9nK�9�I�9�H�9�J�9�I�9gI�9�G�9�I�9�I�9gG�9�I�9rH�9	H�9)J�9�H�9�I�9yJ�9-J�9x   x   �M�9�H�9
G�9�G�9�J�9,K�9J�9K�9	K�9�K�9�H�9~F�9�H�9�L�9&I�9�I�9hI�9�K�9RO�9rH�9%K�9�K�9�J�9XK�9�H�9oN�9VK�9�H�9�I�9�I�9x   x   rJ�9{E�9eK�9J�9L�9PH�9�G�9-H�9TK�99H�9�K�9�E�9_J�9�I�9�G�9zI�9�G�9VO�9�K�9�G�9�M�9�H�9 N�9�H�9�K�9�O�9�H�9%I�9`H�9�H�9x   x   2H�9�L�9[I�9kG�9G�9�K�9�J�9�G�9I�9�I�9;L�9H�9H�9�H�9M�9#H�9�I�9pH�9�G�9P�9�L�9TM�9�N�9G�9DI�9�H�9hH�9�L�9NI�9PH�9x   x   pK�9I�9I�9KK�9�I�9O�9�J�9_I�9lH�9�H�9*L�9J�9�H�9K�9OL�9L�9�I�9&K�9�M�9�L�9�M�9�L�9�O�9�J�9�I�9L�9lL�9�J�9GI�9�I�9x   x   �I�9�E�9I�9�G�9�G�97G�9eH�9]J�9PF�9�I�9�I�9LJ�9�H�9MG�9M�9oI�9gG�9�K�9�H�9UM�9�L�9�G�9�J�9RG�9]J�9�L�9�G�9�H�9�I�9K�9x   x   �H�9=I�9�J�9�F�9bF�9TF�9J�9'H�9�H�9-I�9�F�9�J�9�H�9lJ�9TJ�9�K�9�I�9�J�9�M�9�N�9�O�9�J�9_K�9�J�9�I�9JJ�9�H�9RK�9�F�9�H�9x   x   �F�9M�9-L�9H�9�H�9KL�9�M�9�G�9
G�9�G�9J�9L�9 M�9�I�9�G�9�K�9tH�9\K�9H�9G�9�J�9SG�9�J�9�H�93J�95M�9�K�9bJ�9MG�9�G�9x   x   �I�9 H�9�G�9bH�9�F�9�G�9�H�9�E�9�J�9LI�9BI�9�I�9�J�9+K�9pI�9J�9H�9�H�9�K�9CI�9�I�9[J�9�I�9-J�9�I�9�I�9�H�9�I�9"K�9�E�9x   x   GJ�9�F�9L�9ML�9�G�9aJ�9 K�9`K�9�K�9�G�9�K�9�I�9�K�9�J�9�L�9�L�9'J�9rN�9�O�9�H�9L�9�L�9NJ�93M�9�I�9�L�9�G�9YK�9K�9!K�9x   x   dE�9�H�9zI�9�G�9�D�9I�9=I�9E�9B�9�G�9<I�9�L�9.I�9MG�9�K�98G�9�H�9TK�9�H�9iH�9lL�9�G�9�H�9�K�9�H�9�G�9NB�9�E�9�I�9H�9x   x   �J�9sJ�9�J�9�K�9NG�9PF�9CG�9�E�9IK�9�I�9�H�9�J�9^H�9�K�9�M�9�H�9�I�9�H�9#I�9�L�9�J�9�H�9PK�9aJ�9�I�9UK�9�E�9�E�9�F�9H�9x   x   �G�9�J�9�F�9�H�9�G�9<F�9�H�9�K�9�J�9H�9�G�93J�9/I�9OG�9FI�9�H�9|J�9�I�9aH�9OI�9EI�9�I�9�F�9LG�9%K�9K�9�I�9�F�9xG�9H�9x   x   �J�9L�9�B�9nG�9TH�9�H�9�K�93E�9`G�9H�9J�9�I�9�I�9�H�9�I�9�J�9/J�9�I�9�H�9RH�9�I�9K�9�H�9�G�9�E�9!K�9H�9H�9 H�9�B�9x   x   ��9�9�9t�9X �9��9c�9:$�9!�9�9��9a�9=!�9��9��9�#�9��9k�9- �9� �9"�9��9 �9�"�9��9��9c �9��9|�97�9x   x   �9��9��9-"�9�"�9��9V�9*�9�!�9�9M�9��9X�9N!�9� �9B!�9��9�9��9��9��9>!�9��9U�9��9#�9D"�9��9��9&�9x   x   �9��9
�9f�9��9��9�9#�9i#�9��9�$�9� �9T"�9+$�9��9	%�9�"�9�!�9$�9��9�#�9v!�9��9w �9��9��9:�9I�9@�9� �9x   x   p�9*"�9d�9��9�!�90�9��9��9��95�9!�9��9�!�9� �93�9�!�9 �9� �9N�9(�9��9��9��9j!�9��9��9� �9�9S�9~�9x   x   Z �9�"�9��9�!�9� �9��9��9,�9 �9��9\�9|�9��9Q�9v �9��9.�9�9� �9��9��9 �9@ �9�!�9p�9�#�9( �9��9�$�9��9x   x   ��9��9��90�9��9��9��9� �9W�9��9�!�9<"�9
�9e�9!�9e!�9 �9u�9X!�9��9� �9��9; �9y �9g�9�9��9�9i�9x�9x   x   `�9Z�9�9��9��9��9v�9�!�9��9P"�9"�9U!�9"�9� �9=#�9.!�9:�9[!�9U�9#�9��9��9��9�9��9��9� �9��9��9��9x   x   8$�9&�9#�9��9/�9� �9�!�9.�9v�9*!�9g�9��9�9��9�!�9��9��9�"�9Y!�9P�9��9�#�9J�9$�9s!�9��9�"�9#�9+�9
"�9x   x   !�9�!�9g#�9��9 �9Z�9��9s�9��9�9��9{�9V �9*�9y�9��9��9s�9��9s�9�!�9�!�9��9�#�9��9!�9�$�9:�9��9#�9x   x   �9 �9��90�9��9��9K"�9(!�9�9 �9��9��9I!�9��9u �9�"�9��9��9��9O�9��9 �9��9��9�9�"�9;"�9J�9� �9s�9x   x   ��9H�9�$�9!�9_�9�!�9"�9`�9��9��9��9��9A�9��9"�9!�9��9Q"�9'$�9��9��9� �9� �9"�9��9.�9�9^!�9�!�9� �9x   x   e�9��9� �9��9|�9="�9S!�9��9}�9��9��9^�9B�9!�9Z"�9��91�9#!�9� �9� �9��9R�9��9� �9��9��9H!�9��9��9 �9x   x   >!�9W�9T"�9�!�9��9
�9"�9�9U �9H!�9=�9C�92!�9��9G�9 #�99#�9s�9 �9�"�9� �9I"�9J�9��9��9��9��9�"�9��9l#�9x   x   ��9Q!�9,$�9� �9R�9d�9� �9��9.�9��9��9!�9��99�9 �9#�9[!�9��9�"�9��9�!�9� �9W�9e!�9"�9Q�9# �9:"�9��9"�9x   x   ��9� �9��94�9{ �9~!�9:#�9�!�9y�9v �9"�9]"�9H�9 �9��98!�9��9��9�!�9��9�9�9Q#�9N�9�#�9�9��9�9"�9| �9x   x   �#�9D!�9%�9�!�9��9d!�9-!�9�9��9�"�9!�9��9�"�9#�98!�9$�9��9� �9�#�9�!�9A�9#�9{�9��9/"�9��9#!�9�"�9� �9��9x   x   ��9��9�"�9�9-�9 �98�9��9��9��9��9.�96#�9Z!�9��9��9+ �9�!�9�!�9[!�9"�9� �9#�90"�9�!�9�!�9z"�9�"�9 �9i�9x   x   k�9 �9�!�9� �9�9z�9Y!�9�"�9q�9��9O"�9!!�9t�9��9��9� �9�!�9��9�9`"�9��9
#�9�!�9��99"�9]�9�9� �9�!�9i�9x   x   1 �9��9$�9L�9� �9Z!�9Q�9]!�9��9��9+$�9� �9 �9�"�9�!�9�#�9�!�9�9�$�9 �9��9��9%�98 �98%�9��9�"�9e#�9�!�9�!�9x   x   � �9��9��9*�9��9��9 �9O�9q�9P�9��9� �9�"�9��9��9�!�9[!�9d"�9 �9� �9��9��9? �9��9�!�9N �9�!�9��9q �9�"�9x   x   �9��9�#�9��9��9� �9��9��9�!�9��9��9��9� �9�!�9�9B�9"�9��9��9��9O!�9��9��9��9�#�9��9��9� �9T�9��9x   x   �9C!�9|!�9��9 �9��9��9�#�9�!�9�9� �9R�9H"�9� �9	�9#�9� �9#�9��9��9��9�9h"�9��9(#�9��9]!�9#�9��9]!�9x   x    �9��9��9��9A �9: �9��9Q�9��9��9� �9��9H�9X�9L#�9}�9#�9�!�9$�9> �9��9i"�9�$�9��92$�9��9��9��9w�9 �9x   x   �"�9Y�9z �9j!�9�!�9y �9�9$�9�#�9��9"�9� �9��9j!�9J�9��9/"�9��9: �9��9��9��9��9z�9O!�9��9t �9#�9��9\#�9x   x   ��9��9��9��9r�9j�9��9t!�9��9�9��9��9��9"�9�#�9."�9�!�98"�97%�9�!�9�#�9$#�95$�9K!�9��9��9��9��99�9�"�9x   x   ��9#�9��9��9�#�9�9��9��9�9�"�9*�9��9��9S�9�9��9�!�9d�9��9Q �9��9��9��9��9��9f�9�!�9��9T�9��9x   x   c �9E"�9=�9� �9( �9��9� �9�"�9�$�99"�9�9G!�9��9& �9��9!!�9r"�9�9�"�9�!�9��9[!�9��9t �9��9�!�9%�9�"�9�!�9S�9x   x   ��9��9J�9�9��9�9��9#�9=�9K�9b!�9��9�"�97"�9�9 #�9�"�9� �9f#�9��9� �9	#�9��9
#�9��9��9�"�9��9I�9� �9x   x   y�9��9;�9V�9�$�9g�9��9)�9��9� �9�!�9��9��9��9 "�9� �9
 �9�!�9�!�9n �9P�9��9}�9��96�9Y�9�!�9L�9<$�9u�9x   x   7�9(�9� �9��9��9v�9��9"�9#�9u�9� �9 �9n#�9"�9| �9��9d�9k�9�!�9�"�9��9Y!�9 �9[#�9�"�9��9M�9� �9w�9� �9x   x   ��93��9���9���9��9���9>��9���9��9���9���9���9d��9���9���9��9n��9��9���9��9S��9���9V��94��9��9���9D��9���9���9|��9x   x   +��9���9���9���9i��9Y��9���9l��9���9>��9���9X��9'��9���9d��9���9���9���9���9���9���9h��9���9^��9��9���9���9\��9e��9���9x   x   ���9���9���9���9F��9/��9j��9v��9���9���9���9���9���9\��9^��9���9���9���9���9���9���9��9 ��9w��9w��9���9���9{��9��9��9x   x   ���9���9���9��9���9���9J��9-��9���9���93��9���9W��9F��99��9L��9���9E��9/��9���9��9��9���9��9��9k��9���9|��9���9���9x   x   ��9h��9F��9���9���9���9���9r��9	��9���9'��9���9���9 ��9��9t��9q��9x��9D��9)��9���9[��9���9���9a��9S��9���9"��9���9���9x   x   ���9[��9+��9���9���9!��9���9���9K��9m��9���9i��9h��9B��9���9���9���9��9{��9���9���9x��9���9V��9���9���9���9���9���9���9x   x   :��9���9k��9K��9���9���9��9���9���9���9+��9���9���9d��9���9���9���9v��9���9M��9���9���9���9P��9M��9���9���9��9��9���9x   x   ���9h��9y��93��9o��9���9���9���9��9���9���9���9���9��99��9��9���9~��9���9��9A��9���9��9z��9V��9���9l��9���9���9B��9x   x   ���9���9���9���9��9M��9���9��9���9���9���9g��9+��9���9��9e��9���9o��9 ��9G��9���9���9���9���9��9��9���9���9��9���9x   x    ��9D��9���9���9���9j��9���9���9���94��9q��9���9���97��9���9��9���9���9��9���9���9��9��9���9���9��9��9���9}��9���9x   x   ���9���9���94��9"��9���9,��9���9���9n��9���9P��9���9���9���9���9:��9���9���9k��9���9x��9���9^��9���9j��9i��9���9c��9���9x   x   ���9W��9���9���9���9f��9���9���9d��9���9T��9���9���9���9���9+��9���9���9���9���9���9��9���9J��9���9��9��9R��9R��9���9x   x   f��9)��9���9Y��9���9e��9���9���9/��9���9��9���9!��9	��9���9���9���9���9���9���9Z��9���9s��9���9���9���9`��9j��9Q��9���9x   x   ���9���9Y��9F��9 ��9@��9g��9��9���96��9���9���9��9���9��9f��9���9���9*��9���9F��9A��9Z��9���9i��9���9_��9t��9N��9/��9x   x   ���9c��9^��98��9���9���9���9;��9��9���9���9���9���9��9L��9;��9<��9���9���9!��9���9s��9t��9���9`��9o��9D��9 ��9-��9
��9x   x   ���9���9���9M��9u��9���9���9��9b��9��9���9,��9���9i��9>��9���9���9���9v��9���9���9���9���9���9���9���9,��9'��9���9���9x   x   n��9���9���9���9o��9���9���9���9���9���9>��9���9���9���9:��9���9���9_��9n��9���9���9Y��9��9k��9\��9���9��9(��9��9���9x   x   ��9���9���9H��9y��9��9z��9���9k��9���9���9���9���9���9���9���9a��9���9���98��9���9/��9���9��9���9���9T��9���9���9���9x   x   ���9���9���93��9@��9x��9���9���9!��9��9���9���9���9.��9���9t��9p��9���9���9��9���9���99��9���9v��9O��9���9��9���9���9x   x   ��9���9���9���9'��9���9P��9��9J��9���9j��9���9���9���9 ��9���9���98��9��9���94��9W��9���9���9g��90��9\��9?��9\��9���9x   x   Q��9���9���9��9���9���9���9B��9���9���9���9���9]��9G��9���9���9���9���9���9.��9���9A��9���9!��9]��9���96��9���9���9<��9x   x   ���9e��9���9��9Z��9z��9���9���9���9��9x��9��9���9B��9s��9���9T��9.��9���9Y��9F��9���9���9���9-��9���9���9z��9��9��9x   x   W��9���9��9���9���9��9���9��9���9��9���9���9q��9Z��9q��9���9��9���96��9���9���9���9���9���9���9��9���9���9���9/��9x   x   5��9_��9u��9��9���9U��9O��9{��9���9���9]��9K��9���9���9���9���9k��9��9���9���9!��9���9���9���9H��9���9���9���9@��9?��9x   x   ��9��9t��9��9\��9���9P��9S��9��9���9���9���9���9k��9c��9���9]��9���9w��9f��9`��9.��9���9I��9;��9���9���9���9]��9���9x   x   ���9���9���9m��9V��9���9���9���9��9��9l��9"��9���9���9h��9���9���9���9M��9-��9���9���9��9���9���9���9r��9���9���9���9x   x   E��9���9���9���9���9���9���9m��9���9��9g��9��9^��9`��9D��9)��9��9T��9���9X��95��9���9���9���9���9o��9B��9���9��9���9x   x   ���9[��9u��9w��9!��9���9��9���9���9���9���9R��9k��9{��9#��9)��9*��9���9#��9A��9���9}��9���9���9���9���9���9a��9���9f��9x   x   ���9l��9��9���9���9���9��9���9��9~��9`��9S��9S��9J��9+��9���9��9���9���9[��9���9��9���9>��9]��9���9��9���9���9���9x   x   w��9���9��9���9���9���9���9>��9���9���9���9���9���92��9��9���9���9���9���9 ��9>��9��9/��9@��9��9���9���9c��9���9��9x   x   ���9S��9;��9��9���9���9z��9���9���9���9��9���9��9!��9f��9���9Y��9
��9���9���9���9)��9���9	��9���9���9{��9���9���9���9x   x   V��9���9P��9���9���9���9���9���9��9���9���9��9���9��9%��9N��9w��9Q��9���9���9��9E��9���9���9���9���9L��9���9���9J��9x   x   ;��9O��9���9���9q��9���9(��9_��9k��9*��9
��9���9 ��9V��9<��9D��9��9���9*��9���9+��9^��9���9���9���9S��9v��9L��9���9��9x   x   ��9���9���91��9��9���9���9���9���9D��9���9���9���9���9���9=��9���9A��9��9��9��9~��9���9w��9h��9W��9M��9 ��9l��9V��9x   x   ���9���9o��9"��9���91��9���9���9���9���9���94��9k��9���9t��9-��9z��9���9���9���9��9���9��9��9?��9z��9x��9���9���9t��9x   x   ���9���9���9���91��9���9��9$��9���97��9���9���9���9��9��9��9_��94��9��9���9���9��9+��9y��9���9Z��9F��9���9���9 ��9x   x   |��9���9+��9���9���9
��9|��9"��9��9+��9���9���9��9���9���9���9E��9I��9���9H��9*��9���9q��9���9���9��9���9R��9���9���9x   x   ���9���9]��9���9���9$��9��9���9d��9���9���9Q��9H��9-��9��9���9���9|��9��90��9.��9\��9���9���9���9��9���9���9���9���9x   x   ���9��9g��9���9���9���9��9e��90��9{��9���9���9]��9���9,��9���98��9��9.��9���9��9v��9]��9���9h��91��9^��9���9���9(��9x   x   ���9���9%��9D��9���95��9,��9���9{��9���9��9F��9w��9��9���92��9��9"��9���9���9���9���9���9���9���9z��9���9��9���9���9x   x   ��9���9��9���9���9���9���9���9���9��9��9���9���92��9���9<��9���9"��9���9R��9^��9���9���9A��9���9(��9��9,��9+��9��9x   x   ���9��9���9���99��9���9���9Q��9���9J��9��9���9^��9m��9$��9���9E��9���9��9U��94��9}��9���9y��9��9���9���9���9���9��9x   x   ��9���9���9���9h��9���9��9F��9\��9q��9���9Z��9���9���9#��9���9���9'��9���9���9r��9���9���9���9���9���9���9K��9���9���9x   x    ��9��9Z��9���9���9��9���9,��9���9��91��9m��9���9���9���9���9���9���9���9���9���9���9v��9���9X��9<��9��9��9��9���9x   x   l��9&��9>��9���9q��9��9���9��91��9���9���9#��9%��9���9���9���9���9P��9���9f��9���9���9V��9���9]��9���9��9���9���9��9x   x   ���9L��9D��9=��9+��9��9���9���9���95��9;��9���9���9���9���9���9y��9=��9.��9���9���9���9:��9C��9���9+��9Z��9���9f��9���9x   x   `��9v��9��9���9|��9`��9E��9���97��9��9���9F��9���9���9���9y��94��9���9���9���9_��9���9���9;��9��9���9���95��9���9z��9x   x   ��9O��9���9<��9���91��9F��9~��9
��9��9��9}��9'��9���9Q��9=��9���9���93��9x��9���9���9���9&��9���9��97��9���9���9���9x   x   ���9���9$��9��9���9��9���9��90��9���9���9!��9���9���9���9)��9���92��9L��9��9���9���9{��9V��9Q��9���9z��9��9���9 ��9x   x   ���9���9���9��9���9���9E��9-��9���9���9P��9Z��9���9���9g��9���9���9w��9��9��9���9^��9���9���9���9"��9,��9���9��9���9x   x   ���9��9-��9��9��9���9%��9*��9#��9���9\��93��9u��9���9���9���9_��9���9���9~��9	��9���9���9a��9��9��9s��9���9��9d��9x   x   (��9E��9^��9~��9���9��9���9`��9w��9���9���9z��9���9���9���9���9���9���9���9^��9���9���9��9���9��9���9���9���9O��9%��9x   x   ���9���9 ��9���9��9)��9r��9���9Z��9���9���9���9���9u��9W��9<��9���9���9z��9���9���9��9 ��9���9��9���9���9��9���9Y��9x   x   
��9���9���9~��9��9{��9���9���9���9���9?��9z��9���9���9���9<��9<��9'��9W��9���9b��9���9���9���9���91��9E��9+��9S��9���9x   x   ���9���9���9k��9A��9���9���9���9e��9���9���9���9���9R��9a��9 ��9��9���9V��9���9��9��9	��9���9���9��9���9���9x��9���9x   x   ���9���9O��9U��9x��9Y��9��9��9-��9y��9)��9���9���9<��9���9*��9���9 ��9���9"��9��9���9���9.��9��9���9���9v��9��9���9x   x   x��9J��9w��9N��9x��9C��9���9���9Z��9���9��9���9���9��9��9W��9���98��9}��9.��9u��9���9���9E��9���9���9���9���9���9���9x   x   ���9���9N��9 ��9���9���9L��9���9���9��92��9���9F��9��9���9���94��9���9��9���9���9���9��9/��9���9w��9���9^��9���9���9x   x   ���9���9���9q��9���9���9���9���9���9���9)��9���9���9��9���9h��9���9���9���9��9��9S��9���9Q��9{��9��9���9���9M��9t��9x   x   ���9C��9��9Y��9r��9 ��9���9���9)��9���9	��9���9���9���9��9���9~��9���9 ��9���9b��9&��9Y��9���9���9���9���9���9r��96��9x   x   ߡ�9���9���9��92��9=��9	��9 ��9���9���9���9���9���9R��9��9B��9���9��9`��9H��9t��9��9ި�9���9˪�9��9M��9¥�9���9���9x   x   ���9M��9ʨ�9���9!��9̦�9��9���9X��96��9è�9���9��9)��9i��9ڨ�9���9���9թ�9���9%��9}��9���9q��9@��9��9��9���9���9��9x   x   ���9Ǩ�9,��9b��9���9ͪ�9Ѧ�9ī�9/��9{��9���9B��90��9���9���9���9ժ�9u��9��9s��9���9_��9Ҧ�9+��9d��9��9���9���9׬�9e��9x   x   ��9���9`��9���9Ԫ�9:��9���9���9��9���9���9���9��9���9��9֪�9���9ͬ�9��9b��9a��9g��9u��9C��9��9���9���9g��9���91��9x   x   5��9#��9���9Ԫ�9I��9 ��9=��9V��9O��9ɪ�9���99��9Z��9���9`��9ë�9x��9f��9���9���9���9ȩ�9���9��9���9���9���9Ǧ�9j��9*��9x   x   9��9̦�9Ϫ�9:��9��9۬�9Ѩ�9��9;��9���9���9���9 ��9��9���9���9���9s��9���9i��9;��9��98��9���9��9���9���9��9���9-��9x   x   ��9��9Ҧ�9���9<��9Ө�9���9���9��9Ū�9���9c��9��9]��99��9@��9���9��9Ƨ�9ק�9H��9D��9s��9˨�9��9\��9���9��9���9
��9x   x   ���9���9ë�9���9Q��9��9���9���9b��9���9D��9��9-��9ͨ�9E��9(��9z��9���9r��9���9I��9ث�9\��9/��9b��9��9D��9���9O��9���9x   x   ��9[��95��9��9O��9>��9��9^��9��9���9S��9{��9���9���9I��9��9¦�9}��9��9ب�9e��9��9��9��9���9���9���9S��9���9���9x   x   ���9:��9{��9���9Ū�9���9ƪ�9���9���9ݫ�9���9���9��9���9ީ�9|��98��9��9��90��9-��9��9���9���9���9��9���9$��9ީ�9`��9x   x   ���9Ũ�9���9���9���9���9���9D��9Q��9���9��9���9��9���9���9%��9y��9��9H��9���9ҫ�9׫�9���9���9+��9K��9
��9!��9U��9���9x   x   ���9���9C��9��9;��9���9b��9��9y��9���9���9���9��9L��9d��9t��9R��9[��9ĩ�9ҩ�9J��9���9j��9���9���9���9}��9N��9l��9٪�9x   x   ���9��92��9��9[��9��9��92��9���9��9���9��9��9֨�9M��9T��9���9��9H��9���9���9���9r��9��95��9���9%��9[��9`��9#��9x   x   S��9(��9���9���9���9��9]��9̨�9���9���9���9N��9֨�9Ϋ�9���9ܩ�9i��9:��9���9B��9���9��9$��9��9���98��9Ƭ�9 ��9���9��9x   x   ��9d��9���9��9a��9���98��9A��9I��9٩�9���9a��9N��9���9���9!��9/��9���9��9Ԩ�9]��9Ш�9���9ܪ�97��9���99��9��9Χ�95��9x   x   >��9ب�9���9ت�9ū�9���9>��9&��9��9|��9*��9v��9T��9ک�9%��9��9���9���9���9ͨ�9��9���9��9I��9���9$��9I��99��9��9~��9x   x   ���9���9Ԫ�9���9z��9���9æ�9|��9���94��9|��9T��9���9i��90��9���9��9V��9���9��9���9̪�9Ъ�9���9V��93��9��9/��9l��9���9x   x   ��9���9v��9ͬ�9`��9s��9��9���9}��9��9���9Z��9��98��9��9���9U��9/��9���9#��9U��9���9ٮ�9���9���9��9N��9��9	��9���9x   x   _��9ש�9��9��9���9��9Ƨ�9v��9��9��9L��9©�9E��9���9���9���9{��9���9���9��9M��9��9���9A��9��9���9���9���9��9��9x   x   D��9���9v��9a��9���9k��9ۧ�9���9Ө�92��9���9ө�9©�9@��9ڨ�9Ш�9��9%��9��9��9g��9��9��9Ī�9۩�9e��9 ��9|��9ĥ�9q��9x   x   v��9"��9���9b��9���98��9I��9M��9_��9(��9Ы�9K��9���9���9^��9��9���9T��9Q��9k��9��9`��9���9��9��9���9X��9��9۩�9��9x   x   ��9y��9b��9c��9̩�9��9E��9ܫ�9��9���9ݫ�9���9���9��9Ѩ�9���9̪�9���9��9��9Y��9	��9��9���9;��9���9���98��9ɨ�9��9x   x   ۨ�9���9Ԧ�9q��9���94��9t��9]��9��9���9���9l��9s��9$��9���9��9ת�9֮�9���9��9���9��9��9ɩ�9���9��9���9���9ȩ�9V��9x   x   ���9n��9.��9@��9��9���9ʨ�92��9��9���9���9���9��9��9��9G��9���9���9?��9ª�9��9���9ͩ�9���9C��9��9A��9���9���92��9x   x   Ϊ�9B��9e��9|��9���9��9��9c��9���9���9,��9���97��9���98��9���9T��9���9��9ة�9��9<��9���9F��9���9���9Ԫ�9(��9Ƥ�9K��9x   x    ��9��9��9���9���9���9\��9��9���9��9G��9���9��95��9���9$��94��9��9���9d��9~��9���9��9$��9���9!��93��9��9)��9���9x   x   P��9��9���9���9���9¨�9���9C��9���9���9��9z��9)��9Ǭ�98��9K��9��9L��9���9 ��9U��9���9���9C��9Ԫ�93��9���9`��9Ԫ�9 ��9x   x   ĥ�9���9���9f��9Ȧ�9��9��9���9Q��9&��9#��9J��9X��9���9��98��91��9	��9���9|��9��96��9���9���9%��9��9g��9���9���9���9x   x   ���9���9Ҭ�9���9e��9���9���9L��9���9٩�9T��9p��9d��9���9Ч�9��9m��9��9��9ɥ�9��9ʨ�9Ʃ�9���9���9(��9֪�9���9���9I��9x   x   ��9���9c��93��9+��92��9��9���9���9a��9���9ت�9"��9v��95��9y��9{��9���9��9o��9��9��9U��91��9G��9���9��9���9R��9Q��9x   x   ���9%��9x��9̆�9���9?��9>��9��9ȃ�9���9O��9��9O��9���9�9x��9J��9G��9��9��9���9\��9��9��9҅�9��9��90��9��96��9x   x   #��9��90��9��9ڂ�9��9��9Æ�9n��9��9ކ�9���9��91��9|��9X��9���9Չ�9*��9n��9���9s��9V��9׉�9���9��9-��9���9��9O��9x   x   w��90��9���9*��9���96��9|��9O��94��9��9;��9Ӄ�9��9���9H��9	��9��9�9E��9��9��9���9���9Ӄ�9���9���9u��9m��9��9���9x   x   ͆�9��9,��9|��9H��9��9+��98��9��9���9n��9��9���90��9��9Ճ�93��9;��9���9w��9-��9̈�9���9��9��9���9�9���9(��9΀�9x   x   ���9ق�9���9F��9��9���9ȃ�9Ї�9>��9��9q��9���9r��9\��9܈�9Z��9���9p��9̈́�9g��9��93��9���9���9ʇ�9���9���9��9U��9��9x   x   >��9��94��9|��9���9y��9���9��9���9J��9]��9'��9K��9=��9Ӈ�9���9���9���9G��91��9���95��9���9���9E��9[��9Z��9̈́�9w��9%��9x   x   >��9��9~��9-��9Ƀ�9���9��9ņ�9���92��9ۃ�9F��9Ԅ�9'��9ւ�9@��9���9��9g��92��9ل�9 ��9���9j��9.��9���9���9v��9C��9���9x   x   ��9�9T��99��9Ї�9��9Ć�9���9n��9��9ɇ�9҆�9ц�9���9���9܃�9���9w��9���9���9���9��9P��9��9��9���9���9���9u��9ʄ�9x   x   ˃�9k��9.��9��9=��9���9���9j��9���9���97��9.��9Y��9/��9��9���9���9B��9���9Ƈ�9(��9��9���9h��9���9?��9��9��9l��9͂�9x   x   ��9��9��9���9��9J��94��9��9���9���9R��9���9ڂ�9���9���9Ä�9J��9]��9U��9چ�9���9ք�9Y��9���9U��9>��9��9@��9͆�9���9x   x   N��9ކ�9;��9r��9t��9[��9݃�9ɇ�97��9T��95��9a��9/��9͇�9i��9��9B��9O��9n��9��96��9G��9���9���9��9���96��9��9���9��9x   x   ��9���9σ�9��9���9(��9E��9҆�9.��9���9_��9���9j��9���9���9���9���9ł�9���9��9���9��9Ń�9?��9ه�9@��9F��9���9��9���9x   x   M��9��9��9���9t��9L��9ׄ�9І�9W��9܂�9-��9h��9��9���9��9���9���9��9]��9ӄ�9]��9i��9/��9���9��9���9���9D��9+��9���9x   x   ���93��9���94��9\��99��9'��9���9+��9���9͇�9���9���9F��9Z��9���9���9���98��9z��9W��9���9���9Ӄ�9���9��9���9:��9���9��9x   x   �9���9G��9��9ވ�9ԇ�9܂�9���9��9���9l��9���9���9W��9x��9q��9��9n��9��9���9���9��9���9S��9���9���9���9X��9׈�9_��9x   x   u��9a��9��9Ӄ�9V��9���9@��9܃�9Ä�9Ą�9��9���9���9���9t��9���9��9Z��9��91��9���98��9L��9���9���9��9��9���9#��9~��9x   x   G��9���9
��93��9���9���9���9���9���9H��9@��9���9���9���9��9��9_��9Å�9��9���9҄�9���9=��9��9���9z��9���9Q��9<��9���9x   x   G��9׉�9���9>��9t��9���9��9w��9G��9c��9O��9Ƃ�9��9���9o��9Y��9Ņ�9<��9U��9���9u��9
��9���91��9k��9��9%��9e��9��99��9x   x   ��9&��9A��9��9ʄ�9A��9j��9���9���9R��9i��9���9_��9>��9���9��9��9U��9��9j��9��9���9>��9���9���9*��9���9<��9Շ�9���9x   x   ��9p��9���9y��9c��9-��92��9���9ɇ�9ۆ�9��9��9Մ�9z��9���92��9���9���9g��9I��9h��9���9��9B��9��9���9��9V��9h��9���9x   x   ���9���9��9-��9���9���9؄�9���9,��9���96��9���9a��9W��9���9���9ф�9x��9��9h��9���9S��9���9ˆ�9���9-��9}��9=��9o��9���9x   x   _��9x��9���9ˈ�94��95��9��9߁�9��9ք�9E��9��9k��9���9��9:��9���9��9���9���9R��9���9���9Ɇ�9��9���9��9ۃ�9���9���9x   x   ��9T��9���9Ć�9���9���9���9N��9���9W��9���9�9/��9���9���9K��9>��9���9=��9��9���9���91��9Ƈ�9f��9���9S��9���93��9��9x   x   ��9Չ�9у�9��9��9���9i��9��9h��9���9���9A��9���9Ӄ�9U��9���9��93��9��9D��9Ɇ�9ņ�9Ƈ�9���9݃�9f��9���9V��9��9��9x   x   Յ�9���9���9��9ɇ�9C��90��9��9���9Q��9��9܇�9���9���9���9���9���9m��9���9���9���9��9f��9ރ�9L��9���9\��9^��9L��9���9x   x   ��9��9��9���9���9X��9���9��9B��9<��9���9D��9���9��9���9��9x��9��9+��9���9.��9���9���9c��9���9��9t��9N��9p��9~��9x   x   ��9*��9m��9���9���9R��9���9���9��9��97��9F��9���9���9���9��9���9%��9���9���9���9��9S��9���9[��9u��9���9#��9���9r��9x   x   4��9���9n��9���9��9̄�9x��9���9��9=��9��9���9G��9;��9T��9 ��9R��9e��9;��9W��9=��9݃�9���9V��9_��9L��9!��9΄�9ȅ�9���9x   x   ��9��9��9,��9U��9v��9B��9w��9s��9І�9���9��9*��9���9Ԉ�9"��9;��9��9ԇ�9g��9m��9���96��9$��9S��9m��9���9̅�9���9r��9x   x   5��9K��9���9р�9��9!��9���9ʄ�9΂�9���9��9���9���9��9a��9���9���98��9���9���9���9���9��9��9���9���9r��9���9r��9���9x   x   �f�9c�9ne�9�d�9mc�9|c�9�_�9�`�9�g�96c�9�`�9�b�9�_�9�`�9Qb�9�_�9�a�9T_�9�_�9#b�9�a�9Dc�9�g�9�`�9�`�91d�9�b�9�d�9�c�9�b�9x   x   c�9�`�9ka�9�_�9qc�9f�9�^�9Lc�9�b�9Oa�9�d�96d�9�c�9�a�9	c�9$c�9�b�9�d�9;d�9Ud�9�`�9c�9�b�9�_�9�d�9�b�9W`�9b�9b�9tb�9x   x   ne�9ja�9c�9f`�9�^�9M`�9`�9�d�9b�9�e�9�a�9�b�9�b�9`�9Gb�9@_�9�a�9�a�9c�9f�9b�99e�9�_�9�_�9�`�9�`�9�a�9�`�9�d�9�a�9x   x   �d�9�_�9g`�9Va�9>e�9p`�9�c�9�d�9tc�9�d�9�b�9�e�9d�9a�9�a�9�d�9�f�9ib�9�c�9�c�9d�9nc�9�`�9Ie�9_�9�`�99a�9d�9�c�9�b�9x   x   hc�9nc�9�^�9Ce�9�g�9�a�9�c�9h`�95b�9Ic�98b�9]a�9�`�9�^�9�_�9�`�9b�9'd�9gb�9�`�98d�9Sa�9�g�9�e�9�`�9b�9�b�9d�9�e�9�c�9x   x   �c�9f�9M`�9s`�9�a�9ia�9�b�9�b�9�d�9�a�9�b�9Cd�9Jd�9�d�98e�9�b�9a�9!e�9�a�9Mb�9sa�9�a�9o`�9�_�9e�9|d�9k`�9�_�9a�9�_�9x   x   �_�9�^�9`�9�c�9�c�9�b�9c�9�a�9�c�9�c�9@g�9a�9�_�9�`�9zf�9	e�9ic�9�a�9d�9�b�9�c�9�c�9)`�9�^�9	a�9ba�9�a�9�c�9q`�9c�9x   x   �`�9Jc�9�d�9�d�9j`�9�b�9�a�9�^�9�`�9vb�9Ba�9'b�9�a�9�a�9�a�9t`�94_�9a�9Fb�9>`�9�d�9d�9�c�9C`�9�b�9�^�9�b�9
c�9�^�9Yc�9x   x   �g�9�b�9b�9rc�95b�9�d�9�c�9�`�9�a�9la�9tc�9�c�9Mc�9Ib�9�a�9�`�9�c�9,e�9�b�9rc�9�b�9�b�9�g�9&d�9�b�9�`�9(c�9b�9�`�9yd�9x   x   5c�9Ua�9�e�9�d�9Ic�9�a�9�c�9rb�9ha�9je�9�e�9�f�9d�9�`�9�b�9bc�9�a�9�b�9�d�9e�9sa�9�b�9of�9"_�9Q_�9�c�9�a�9j`�9�`�9[e�9x   x   �`�9 e�9�a�9�b�9:b�9�b�9;g�9Ba�9vc�9�e�9�h�9�e�9�d�9�`�9fg�9�b�9Jb�9�b�9�b�9e�9�`�9�`�9�b�9Db�9(b�9d�9�b�9�`�9Bb�9�a�9x   x   �b�98d�9�b�9�e�9\a�9Gd�9a�9'b�9�c�9�f�9�e�9@c�9Sa�9�`�9kd�9�`�9'f�9�a�9�c�9/b�9�c�9�c�9*c�9�c�9Y_�99`�9�c�9d�9bd�9�b�9x   x   �_�9�c�9�b�9d�9�`�9Ld�9�_�9�a�9Oc�9d�9�d�9Pa�9�`�9�c�9Xa�9�c�9�b�9�c�9�`�9�c�9e�9�d�9�b�9c�9``�94b�9jc�9Wc�9%e�9fd�9x   x   �`�9�a�9`�9a�9�^�9�d�9�`�9�a�9Jb�9�`�9�`�9�`�9�c�9�^�99a�9�_�9�a�9�_�9]`�9Id�98]�9=a�9�b�9�d�9�d�9�b�9Wa�9b^�9�c�9�_�9x   x   Vb�9	c�9Db�9�a�9�_�99e�9tf�9�a�9�a�9�b�9cg�9jd�9Za�96a�9�b�9�b�9�b�9�`�98b�9�d�9�a�9�e�9�a�9�a�9�a�9=e�9�a�9tc�9�b�9�`�9x   x   �_�9!c�9>_�9�d�9�`�9�b�9e�9u`�9�`�9ac�9�b�9�`�9�c�9�_�9�b�9A_�9Mb�9�d�9	c�9d�9]c�9'b�9Ha�9�`�9�b�9�c�9id�9 d�9�c�9(b�9x   x   �a�9�b�9�a�9�f�9b�9a�9ic�93_�9�c�9�a�9Ib�9'f�9�b�9�a�9�b�9Nb�9�d�9c�94a�9�a�9b�9Kf�9g�9�e�9�a�9Ga�9{`�9�b�9f�9/b�9x   x   V_�9�d�9�a�9ib�9&d�9 e�9�a�9a�9,e�9�b�9�b�9b�9�c�9�_�9�`�9�d�9c�9b�9kb�9<c�9e�9b�9c�9Te�9�c�9
c�9b�9c�9|c�9�a�9x   x   �_�9>d�9c�9�c�9lb�9�a�9d�9Db�9�b�9�d�9�b�9�c�9�`�9Z`�98b�9	c�97a�9lb�9�`�9Nc�9�b�9Wc�9�a�9c�9�_�9>b�9�`�9�c�9�b�9^`�9x   x   %b�9Yd�9f�9�c�9�`�9Ob�9�b�9=`�9wc�9e�9e�90b�9�c�9Gd�9�d�9d�9�a�9<c�9Mc�9�`�9�c�9�c�9�a�9�c�9�c�9�a�9d�9ud�9�b�94e�9x   x   �a�9�`�9b�9d�9:d�9ua�9�c�9�d�9�b�9ma�9�`�9�c�9e�9=]�9�a�9_c�9b�9"e�9�b�9�c�9`�9tc�9
a�9$e�9za�9�c�9Ua�9�^�9�d�9�b�9x   x   >c�9c�98e�9nc�9Oa�9�a�9�c�9d�9�b�9�b�9�`�9�c�9�d�9;a�9�e�9(b�9Gf�9b�9Wc�9�c�9wc�98d�9�b�9�f�9Yb�9yf�9c`�9d�9�c�9�`�9x   x   �g�9b�9�_�9�`�9�g�9k`�9+`�9�c�9�g�9mf�9�b�9+c�9�b�9�b�9�a�9La�9g�9c�9�a�9�a�9a�9�b�9�e�9ja�9u`�9�c�9c�9?d�9Jc�95e�9x   x   �`�9�_�9�_�9Oe�9�e�9�_�9�^�9B`�9)d�9&_�9Fb�9�c�9
c�9�d�9�a�9�`�9�e�9Ue�9c�9�c�9e�9�f�9fa�9�b�9�d�9xb�9Zc�9V`�9&`�9�d�9x   x   �`�9�d�9�`�9_�9�`�9e�9a�9�b�9�b�9P_�9(b�9V_�9``�9�d�9�a�9�b�9�a�9�c�9�_�9�c�9{a�9Xb�9t`�9�d�9`�9B`�9�c�9�_�9�a�9�a�9x   x   3d�9�b�9�`�9�`�9
b�9zd�9ga�9�^�9�`�9�c�9d�96`�94b�9�b�9=e�9�c�9Ea�9c�9:b�9�a�9�c�9|f�9�c�9vb�9B`�9�a�9c�9`�9�`�9wb�9x   x   �b�9V`�9�a�99a�9�b�9j`�9�a�9�b�9)c�9�a�9�b�9�c�9gc�9Ua�9�a�9jd�9|`�9�b�9�`�9d�9Ra�9c`�9c�9Yc�9�c�9c�9d�9�b�9o_�9n`�9x   x   �d�9b�9�`�9d�9d�9�_�9�c�9c�9b�9h`�9�`�9d�9Uc�9d^�9tc�9#d�9�b�9c�9�c�9td�9�^�9d�9Dd�9W`�9�_�9`�9�b�9�d�9�`�9�c�9x   x   �c�9b�9�d�9�c�9�e�9a�9u`�9�^�9�`�9�`�9Bb�9bd�9"e�9�c�9�b�9�c�9f�9�c�9�b�9�b�9�d�9�c�9Fc�9`�9�a�9�`�9o_�9�`�9�d�9�c�9x   x   �b�9ob�9�a�9�b�9�c�9�_�9c�9Xc�9ud�9Ze�9�a�9�b�9cd�9�_�9�`�9+b�9.b�9�a�9d`�97e�9�b�9�`�95e�9�d�9�a�9ub�9j`�9�c�9�c�9]b�9x   x   )<�9S>�9�B�9Q<�9dA�9=?�9�?�9�B�9R;�9�@�9�E�9O@�9�C�9 E�9lD�9�E�9�C�9�D�9�C�9g?�9F�9�?�9�;�9ZC�9>A�9�?�9�@�9�<�9�@�9>�9x   x   T>�9:D�98?�9SA�9�C�9@�9�B�9�?�9�=�9A�9O=�9�@�9�>�9c>�9SA�9�A�9H?�9?�9{@�9;=�9�A�9S>�9�=�9lB�9�>�9_C�9�A�9�@�9�E�9=�9x   x   �B�95?�9pB�9�C�9X?�9GF�9�@�9dA�9�B�9B<�9�A�9�A�9s?�9TC�9>�9�B�9�>�9yA�9�B�9�;�9B�9XB�9B�9�E�9e@�9�D�9�@�9+>�9WC�9m@�9x   x   S<�9WA�9�C�9�=�9�@�9�@�9=�9UB�9�<�9�?�9�A�9 >�9�C�9C�9\C�9�D�9�>�9�@�9�?�9(>�9�A�9'<�9@�9=A�9�;�9�D�9mC�9i;�9@�9C?�9x   x   eA�9�C�9V?�9�@�9M?�9�?�9B�9�?�9�A�9?�9%@�9A�9|?�9?D�9?�9m@�96@�9�?�9�@�9"@�9C�9�?�9?�9�@�9y@�9�A�9pA�9R<�9)?�9�<�9x   x   <?�9@�9EF�9�@�9�?�9�B�9v?�9C�99B�9�>�9�E�9�=�9*C�9DC�9->�9�E�9!>�9�B�9C�9Z>�9�B�9`@�9�?�9"F�9@�9�?�9B�9�@�9QA�9DA�9x   x   �?�9�B�9�@�9=�9"B�9t?�9F@�94@�9�>�9>�9U?�9�<�9'D�9�<�9�>�9�>�9�=�9?@�9A�9{@�9RA�9 =�9vA�9jA�9oA�9�B�91B�9�B�9B�9<D�9x   x   �B�9�?�9aA�9UB�9�?�9C�92@�9hD�9E�9�?�9@�9SD�9CD�9Q@�9i?�9�E�9�D�9g?�91B�9�?�9�B�9�@�9x@�9B�9�C�9U@�9�@�9A�9[?�9vD�9x   x   Q;�9�=�9�B�9�<�9�A�9<B�9�>�9E�9�D�9�@�9Q@�9{?�9%@�9�A�9]D�9�D�9�>�9BC�9�A�9�<�9C�9=�9�;�9y?�9�?�9�A�9A�9�B�9?�9�?�9x   x   �@�9A�9A<�9�?�9?�9�>�9>�9�?�9�@�9
A�9=�9�=�9&@�9�@�9�@�9�=�9�=�9�>�9h@�9;�9sB�9H@�9�@�9�A�9�A�9`@�9�>�9C�9aB�9�@�9x   x   �E�9K=�9�A�9�A�9"@�9�E�9U?�9@�9O@�9	=�9�:�9=�9�@�9�?�9?�9�F�9�@�9�@�9�B�9Q=�9;E�9R@�9�@�9DC�9	C�9�B�9*C�9B�9�@�9�@�9x   x   M@�9�@�9�A�9�=�9A�9�=�9�<�9TD�9z?�9�=�9=�9}?�9�C�9�=�9�<�9�?�9�>�9�A�9�@�9�?�9�?�9:>�9b>�9�@�9�A�9�B�9�@�9}?�9$>�9Y>�9x   x   |C�9�>�9s?�9�C�9y?�9*C�9'D�9FD�9$@�9#@�9�@�9�C�9XD�9C�9�@�9�C�9P?�9J>�9D�9�?�9v>�9�C�9a>�9�A�9�C�9@�9y>�9�B�9@�9�?�9x   x   �D�9`>�9YC�9C�9=D�9DC�9�<�9X@�9�A�9�@�9�?�9�=�9C�9C�9C�9"C�9?�9%E�96E�9�?�9�C�9[D�9'>�9�@�9�A�9D?�9�D�9�C�9?�9tE�9x   x   jD�9SA�9>�9ZC�9?�9+>�9�>�9g?�9ZD�9�@�9?�9�<�9�@�9C�9�>�9 A�9	D�9�@�9�<�9e@�9z@�9�B�9ZB�9hA�9�A�9A�9aA�9l?�94=�97A�9x   x   �E�9�A�9�B�9�D�9n@�9�E�9�>�9�E�9�D�9�=�9�F�9�?�9�C�9"C�9A�9�E�9o@�9bA�9�C�9�?�9A>�9~@�9�@�9�@�9"B�9U>�9�?�9>E�9�?�9�?�9x   x   �C�9H?�9�>�9�>�96@�9 >�9�=�9�D�9�>�9�=�9�@�9�>�9N?�9?�9D�9o@�9�<�9PA�9�B�9D�9uA�9?>�9�@�9�=�9�@�9�C�9�A�9A�9�>�9�@�9x   x   �D�9?�9wA�9�@�9�?�9�B�9<@�9g?�9@C�9�>�9�@�9�A�9L>�9&E�9�@�9bA�9MA�9�>�9�B�9�@�96>�9	A�9�A�9�=�9B�9�C�9�>�9A�9U?�9�A�9x   x   �C�9y@�9�B�9�?�9�@�9C�9A�92B�9�A�9h@�9�B�9�@�9D�96E�9�<�9�C�9�B�9�B�9c@�9@B�9�A�9�@�9tA�92B�9[>�9rB�9�B�9�D�9�=�9�D�9x   x   d?�97=�9�;�9#>�9!@�9Y>�9z@�9�?�9�<�9";�9Q=�9�?�9�?�9�?�9d@�9�?�9 D�9�@�9BB�9iC�9"A�9�@�9�C�9!C�94B�9D�9�>�9@�9H>�9�@�9x   x   F�9�A�9B�9�A�9C�9�B�9PA�9�B�9C�9tB�9:E�9�?�9t>�9�C�9z@�9A>�9wA�93>�9�A�9#A�9E�9A�9]@�9 >�9�?�9??�9�@�9�D�9?�9?�9x   x   �?�9S>�9XB�9)<�9@�9e@�9 =�9�@�9=�9O@�9R@�99>�9�C�9]D�9�B�9y@�9?>�9A�9�@�9�@�9A�9�A�9�A�9�>�9/A�9�A�9�C�9�C�9�=�9Z@�9x   x   �;�9�=�9B�9@�9?�9�?�9qA�9s@�9�;�9�@�9�@�9c>�9b>�9(>�9[B�9�@�9�@�9�A�9uA�9�C�9\@�9�A�9�?�9�@�9nA�9??�9p>�9/?�9�A�9�@�9x   x   YC�9jB�9�E�9=A�9�@�9$F�9hA�9B�9{?�9�A�9BC�9�@�9�A�9�@�9gA�9�@�9�=�9�=�94B�9%C�9�=�9�>�9�@�9�A�9A�9�@�9o@�9�A�9�A�9�?�9x   x   ;A�9�>�9f@�9�;�9|@�9@�9kA�9�C�9�?�9�A�9	C�9�A�9�C�9�A�9�A�9"B�9�@�9B�9Z>�99B�9�?�91A�9kA�9}A�9C�9C�9�C�9�B�9�@�9�B�9x   x   �?�9^C�9�D�9�D�9�A�9�?�9�B�9R@�9�A�9`@�9�B�9�B�9@�9F?�9A�9T>�9�C�9�C�9nB�9D�9??�9�A�9>?�9�@�9 C�9�@�96@�9@�9[A�9CC�9x   x   �@�9�A�9�@�9nC�9pA�9B�90B�9�@�9A�9�>�9+C�9�@�9x>�9�D�9bA�9�?�9�A�9�>�9�B�9�>�9�@�9�C�9o>�9o@�9�C�94@�9	B�9A�9<A�9 B�9x   x   �<�9�@�9(>�9i;�9V<�9�@�9�B�9A�9�B�9C�9B�9}?�9�B�9�C�9m?�9=E�9 A�9A�9�D�9!@�9�D�9�C�9-?�9�A�9�B�9@�9!A�9�B�9qA�9m<�9x   x   �@�9�E�9VC�9@�9*?�9MA�9B�9W?�9?�9dB�9�@�9%>�9	@�9?�94=�9�?�9�>�9X?�9�=�9G>�9?�9�=�9�A�9�A�9�@�9[A�9=A�9oA�9>�9�?�9x   x   #>�9=�9q@�9F?�9�<�9FA�9;D�9uD�9�?�9�@�9�@�9Y>�9�?�9qE�96A�9�?�9�@�9�A�9�D�9�@�9?�9V@�9�@�9�?�9�B�9FC�9B�9k<�9�?�9B�9x   x   �)�9�!�9��9�"�9s!�9��9 �9V!�9�!�9j �9��9�!�9�9��9c�9^�9��9T�9q�9� �9@�9�9�"�9�"�9< �9��9� �9�#�9��9�!�9x   x   �!�9�9�!�9��9��9�9v�9e#�9�"�9�!�9R�9/ �9�!�9�!�9S�9��9T"�9� �9� �97 �9�"�9�"�9.!�9��9'�9M�9i�9�"�99�9� �9x   x   ��9�!�9v�9`�9!�96�9� �9��9� �9B$�9�!�9� �9�"�9L"�9d �9G"�9#�9u!�9]!�9�"�9W �9��9a"�99�9= �9��9��9� �9�9�9x   x   �"�9��9]�9�&�9��9q#�9�!�9S�9m"�9	!�9� �9��9��9=�9�9y�9��9��9�"�9�#�9p�9� �9)"�9�9�%�9��9;!�9�"�9�!�9v!�9x   x   t!�9��9!�9��9Z�9�"�9r�9�"�9;!�9$ �9�!�9�!�9� �9��9x!�97!�9�!�9� �9��9�"�9� �9�#�9 �9�9/!�9�9�!�9h#�9,"�9�#�9x   x   ��9�96�9n#�9�"�9$�9��9}�9,�9$�9[�9"�9p�9��97"�9��9�#�9��9��9��9��9�#�9w"�9��9y�9��9x!�9)!�9� �9D!�9x   x    �9v�9� �9�!�9r�9��9�"�9��9�!�9� �9� �9�#�9|�9�#�9H �9� �9F!�9��9�!�9�!�9��9[!�9"�9��9. �9�9�9�9m�9��9x   x   W!�9c#�9��9Q�9�"�9�9��9c �9+�9� �9�$�9��9R�9%�9� �9��9n �9��9(�9�"�9��9��9�#�9�!�9G�9�!�9�9v�9� �9L�9x   x   �!�9�"�9� �9p"�9<!�9+�9�!�9%�9��9H �9�9]�9\�9� �9��9��9'"�9��9��97"�9�!�9�!�9 "�9��9� �9@#�9W�9N#�9)!�9��9x   x   j �9�!�9A$�9
!�9% �9
$�9� �9� �9F �9q �9%�9�%�9� �9� �9r!�9� �9�!�9# �9#�9�"�9�"�9� �9 �9�!�9��9F�9��9F �9� �9� �9x   x   ��9S�9�!�9� �9�!�9Z�9� �9�$�9�9%�9t#�9%�9��9`$�9��9 �9
#�9��9�!�9x�9��9��9� �9��9�95�9�9H�9� �9I�9x   x   �!�91 �9� �9��9�!�9"�9�#�9��9`�9�%�9%�9��9M�94%�9!�9��9��9!�9%!�9�!�9*#�9J$�9w!�9 �9��9r�9' �9="�9�#�9�"�9x   x   �9�!�9�"�9��9� �9p�9{�9N�9Y�9� �9��9L�9��9��9#�9^�9�"�9� �9 �9A�9h�9��9^"�9�#�96�9�"�9"�9��9� �9~�9x   x   ��9"�9I"�9;�9��9��9�#�9%�9� �9� �9^$�93%�9��9��9�9"�9�"�9�9��9�"�9X �9��9� �9+�9��9�!�9R�9��9�"�9��9x   x   `�9W�9_ �9�9~!�96"�9K �9� �9��9w!�9��9!�9#�9�9!�9�9�9O �91!�9�!�9� �9L�9�!�9d �9� �9��9�!�9N!�9�!�9� �9x   x   ^�9��9E"�9y�99!�9��9� �9��9��9� �9 �9��9_�9"�9�9��9P!�9)#�97�9��9B!�9� �9�"�9}"�9�"�9�!�9��9��9"�9� �9x   x   ��9U"�9	#�9��9�!�9�#�9C!�9l �9%"�9�!�9#�9��9�"�9�"�9�9P!�9+ �9� �9 �9��9�$�9� �9��9V �9#�9 �98�9� �9r!�9�!�9x   x   T�9� �9u!�9��9� �9��9��9��9��9( �9��9!�9� �9
�9P �9*#�9� �9�"�9��9��9z!�9�!�9y"�9h!�9D�9 �9d"�9� �9G!�9� �9x   x   o�9� �9Y!�9�"�9��9��9�!�9(�9��9 #�9�!�9&!�9�9��9.!�99�9�9��9
#�9��9�!�9B �9D!�9��9�!�9_�9K�9%�9/"�9X�9x   x   � �97 �9�"�9�#�9�"�9��9�!�9�"�93"�9�"�9x�9�!�9@�9�"�9�!�9��9��9��9��9��9��9��9D�9��9��9��9��9�!�9J"�9��9x   x   B�9�"�9X �9t�9� �9��9��9�9�!�9�"�9��9)#�9l�9Y �9� �9A!�9�$�9w!�9�!�9��9�!�9x�9`!�93!�9�"�9�"�9�!�9  �9� �9#�9x   x   �9�"�9��9� �9�#�9�#�9U!�9��9�!�9� �9��9J$�9��9��9P�9� �9 !�9�!�9A �9��9v�9� �9"�9�!�9�!�9��9��9��9r#�9
 �9x   x   �"�91!�9b"�9("�9"�9|"�9"�9�#�9"�9 �9� �9x!�9^"�9� �9�!�9�"�9��9x"�9G!�9D�9`!�9"�9��9�"�9�!�9�!�9�"�9�!�9� �9� �9x   x   �"�9��9;�9�9�9��9��9�!�9��9�!�9��9 �9�#�9(�9i �9z"�9V �9f!�9��9��92!�9�!�9�"�9��9��9:"�9B �9��96 �9��9x   x   ? �9'�9? �9�%�9/!�9|�9, �9J�9� �9��9�9��95�9��9� �9�"�9#�9E�9�!�9��9�"�9�!�9�!�9��9��9��9A�9� �9Z"�9%�9x   x   ��9J�9��9��9�9��9�9�!�9@#�9D�94�9s�9}"�9�!�9��9�!�9�9 �9`�9��9�"�9��9�!�98"�9��9��9\�95!�9"�9l�9x   x   � �9g�9��9=!�9�!�9u!�9�9�9T�9��9�9* �9"�9U�9�!�9��98�9b"�9I�9��9�!�9��9�"�9A �9A�9[�9� �9y�9��9�!�9x   x   �#�9�"�9� �9�"�9d#�9+!�9 �9t�9L#�9D �9F�9<"�9��9��9K!�9��9� �9� �9$�9�!�9 �9��9�!�9��9� �94!�9v�9�9!�9�#�9x   x   ��99�9�9�!�9*"�9� �9k�9� �9)!�9� �9� �9�#�9� �9�"�9�!�9"�9t!�9F!�91"�9I"�9� �9r#�9� �94 �9]"�9"�9��9!�9�!�9�!�9x   x   �!�9� �9}�9x!�9�#�9D!�9��9O�9��9� �9N�9�"�9|�9��9� �9� �9�!�9� �9Z�9��9#�9 �9� �9��9$�9k�9�!�9�#�9�!�9� �9x   x   2��9� �9��9���97��9�9��9:��9@�9D�9%��9�9��9�9��9g�9��9��9��9n�9���9�9��9���9��9�9|��9� �9� �9� �9x   x   � �9 �91�9[�9�9f�9<��9���9���9���9��9�9$�9G�9	�9=�9��9� �9��9��9>��9���9 ��9���9v�9�9�9x�9�9� �9x   x   ��95�9b�9! �9��97��9���9n�9���9+�9;��9j��9� �9���9b�9���95�9h��9��9 �9
��9B�9���9X��9� �9k �9�9~�9+�9��9x   x   ���9[�9 �9 �9��9�9��9��9���9���9	�9J�9���9��9��9g��9@�9< �9���9� �9x�9�9[�9��9� �9���9/�9� �9���94��9x   x   8��9�9��9��94�9���9 �9O�9�9z�99 �9��9��9��9|�9{�9a �9��9���91�9C�9*��9��9��9��9��9���9��9���9���9x   x   �9d�9;��9�9���9[ �9��9���9��9� �9T��9)�9,�9J �9�9���9� �95�9� �9�9���9���9��9��9��9��9��9���9���9]��9x   x   ��99��9���9��9 �9~�9�9.�9|�9��9j��9�9�9l�9B��9��9D�9��9n�9��9���9"�9 �9���9��9v�9|�9O�9��9� �9x   x   8��9���9q�9��9Q�9���92�9z��95�9��9��9� �9� �9���93�9��9���9q�9���9p�9��9��9���9F��9��9�9��9��9$�9��9x   x   9�9���9���9���9�9��9�93�9��9��9� �9f�9, �9�9��9��9s�9!�9V �93��9��9V��9��9�9 �9���9��9���9� �9~�9x   x   E�9���9-�9���9y�9� �9��9��9��93 �9��9��9� �93�9��9��9���9��92 �9� �9���9��9~�9��9M��9�9��9���9 �9�9x   x   #��9��98��9�96 �9Q��9l��9��9� �9��9N��9��9 �9���9���9 ��9N�9 ��9���9Y�9e��9, �9��9}�9*�9��9b�9�9���9h��9x   x   �9�9i��9L�9��9+�9�9� �9e�9��9��9]�9@�9��9X�9� �9W�9��9�9O�9���9=�9�9��9��9C�9w�9��9�9d �9x   x   ��9!�9� �9���9��9*�9�9� �90 �9� �9 �9A�9���99�9w�9���9i �9A�9�9��9��9H �9��9 ��9��9��9��9. �9/�9� �9x   x   
�9D�9���9��9��9F �9o�9���9�90�9���9��97�9E �9��9���9��9��9x��9�9���9��9��9��9M�9��9�90��9i�9���9x   x   ��9�9d�9��9y�9�9C��92�9��9��9���9Y�9w�9��9��9��9��9�9f�99��9n�9��9y�9k �9��9��9��9h��9v�9�9x   x   i�9=�9���9f��9z�9���9��9��9��9��9��9� �9���9���9��9(�9��9� �9� �9D�9��9���9U��9���9��9-�9��9, �9� �9v�9x   x   ��9��96�9C�9` �9� �9E�9���9q�9���9P�9Y�9g �9��9��9��9? �9� �9��9h �9 �9��9q�9�9g��9) �9��9� �9� �9��9x   x   ��9� �9i��97 �9��92�9��9q�9 �9��9��9��9?�9��9�9� �9� �9��9b �9u �9:�9��91 �9��9� �90 �9��9� �9���9��9x   x   ��9��9��9���9���9� �9m�9���9U �94 �9���9�9
�9}��9b�9� �9��9a �9��9� �9�9 �9��9� �9��9���9G�92�9��9U��9x   x   o�9��9 �9� �90�9�9��9n�94��9� �9Y�9R�9��9�9<��9F�9g �9x �9� �9z�9&�9��9�9  �9b�9s �9��96��9��9� �9x   x   ���9A��9	��9v�9E�9���9���9��9���9���9i��9���9��9���9n�9��9  �94�9�9'�9� �9 �9�9��9���9��9e�9���9��9G �9x   x   �9���9B�9�9)��9���9!�9��9V��9��9+ �9>�9D �9�9��9���9��9��9 �9��9 �9���9���9n�9r��9?�9	�97 �9��9G �9x   x   ��9���9���9_�9��9��9 �9���9��9�9��9�9��9��9z�9S��9p�90 �9��9�9�9���9��9���9��9��9��9��9��9��9x   x   ���9���9X��9��9��9��9���9G��9��9��9y�9��9$��9��9m �9���9 �9��9� �9 �9��9s�9���9��9��9l��9�9B�9 �9
�9x   x   ��9q�9� �9� �9��9��9��9��9 �9M��9)�9��9��9P�9��9{��9i��9� �9��9^�9 ��9o��9��9��9	�9��9��9 �9��9� �9x   x   �9�9l �9���9��9��9t�9�9���9#�9��9?�9��9��9��9+�9% �90 �9 �9q �9��9=�9��9k��9��9��9��9���9&�9B�9x   x   ~��9�9�9/�9���9��9{�9��9��9��9c�9y�9��9�9��9��9��9��9J�9��9e�9	�9��9�9��9��9��9�9��9;��9x   x   � �9y�9{�9� �9��9���9O�9��9���9���9�9��9/ �92��9i��9- �9� �9� �97�95��9���98 �9��9H�9 �9���9��9r�9���9���9x   x   � �9�9)�9���9���9���9��9%�9� �9 �9���9�9/�9n�9u�9� �9� �9���9��9��9��9��9��9 �9��9)�9��9���9z��9���9x   x   � �9� �9�91��9���9\��9� �9��9}�9�9i��9h �9� �9���9�9u�9��9��9R��9� �9G �9F �9��9�9� �9B�9:��9���9���9��9x   x   \��9���9]��9^��9���9���9'��9^��9#��9S��9���9;��9R��9��9���9X��9u��9���9���9���9���9��9���9���9	��9)��9���9%��9���9���9x   x   ���9"��9���9���9���9���9���9��9���9���9���9H��9k��9[��9/��9���9%��9���9��9��9<��9���9���9l��9!��9���9 ��9���9���9<��9x   x   _��9���9��9���9��9Z��9(��9��9P��9#��9=��9���9���9B��9#��9���9��9���9U��9X��9+��9���9���9��9���9��9f��9���9��9_��9x   x   Y��9���9���9y��9j��9���9n��9a��9���9��9���9<��9@��9��9C��9p��9���9���9���9���9���9=��91��9���98��9���98��9e��9���9���9x   x   ���9���9��9f��95��9���9?��9���9B��9���9���9��9��9R��9��9���9���9��9D��9���9���9E��9X��9s��9��9���9B��9���9&��9#��9x   x   ���9���9Y��9���9���9���9��9Z��9���9%��9���9���9��9���9���9���9\��9���98��9���9A��9c��9���9���9��9���9���9F��9;��9���9x   x   %��9���9#��9l��9C��9��9K��9���9���9���9��9w��9���9��9
��9]��9���9���9���9z��9���9��9��9m��9���9;��9C��9F��9z��9?��9x   x   d��9	��9��9b��9���9X��9���9���9T��9���9���9+��9���96��9���9���9D��94��9d��9P��9|��92��9���9��9u��9U��9���9���9��9C��9x   x   !��9���9M��9���9D��9���9���9T��9G��9���9���9���9r��9���9��9���9���9
��9N��9���9`��9��9���9B��9���9P��9���9���9>��9���9x   x   T��9���9"��9	��9���9$��9���9���9���9`��9P��9���9��9���9��9��9y��9v��9��9���9���9x��9���9���9k��9x��9M��9���9g��9���9x   x   ���9���9>��9���9���9���9��9���9���9P��9���9a��9��9a��9���9 ��9���9X��9���9���9m��9���9���9���9h��9E��9���9���9���9)��9x   x   =��9H��9���9;��9��9���9s��9)��9��9���9f��9-��9��9���9���9/��9\��9&��9���9��9I��9���9���9q��9���9F��9���9L��9���9���9x   x   R��9j��9���9<��9��9��9���9���9q��9��9��9��9���9���9z��9T��9���9(��9L��9���9h��9���9���9Q��9���9���9���9���9f��9���9x   x   ��9Z��9F��9��9T��9���9��98��9���9���9c��9���9���9��95��9���93��9���9���9I��9d��9��9���9���9���9'��9W��9'��9���9���9x   x   ���9-��9&��9B��9��9���9��9���9���9��9���9���9y��96��9Y��9_��9'��9m��9���9���9���9C��9���9U��9?��9���9M��9���9���9��9x   x   [��9���9���9p��9���9���9Z��9���9���9��9��9-��9U��9���9\��9���9���9���9���9��9E��9���9���9��9��9���9f��9;��9.��9���9x   x   u��9'��9��9���9���9^��9���9F��9���9~��9���9[��9���97��9$��9���9?��9���9p��9���9��9���9���9���9���9���9���9���9���9��9x   x   ���9���9���9���9��9���9���90��9��9p��9W��9!��9&��9���9h��9���9���9%��9���9���9���9���9.��9���9��9���9��98��9v��9��9x   x   ���9��9Z��9���9G��9<��9���9m��9O��9��9���9���9O��9���9���9���9q��9���9���9[��9���9z��9@��9���9���9t��9���9���9��9���9x   x   ���9��9T��9���9���9���9w��9Q��9���9���9���9
��9���9L��9���9��9���9���9[��96��9��9N��9i��9���9���9Q��9��9��9y��9���9x   x   ���9=��9)��9���9���9?��9���9y��9c��9���9k��9I��9d��9c��9���9H��9��9���9���9��9���9)��9��9L��9���93��9���9���9,��9��9x   x   ��9���9���9>��9E��9d��9��93��9��9{��9���9���9���9��9C��9���9���9���9z��9L��9+��9���9A��9���9���9��9���9���9���9���9x   x   ���9���9���9/��9T��9���9 ��9���9���9���9���9���9���9���9���9���9���9+��9>��9f��9
��9<��9��9���9���9o��9���9���9&��9���9x   x   ���9q��9��9���9w��9���9p��9��9B��9���9���9p��9O��9���9O��9��9���9���9���9���9I��9���9���9F��9 ��9���9+��9��9���9���9x   x   ��9&��9���95��9%��9��9���9x��9���9l��9m��9���9���9���9;��9��9���9��9���9���9���9���9���9���9���9D��9���9���9���9���9x   x   #��9���9��9���9���9���99��9T��9O��9s��9H��9H��9���9,��9���9���9���9���9t��9S��94��9��9q��9���9F��9���93��9���9��9o��9x   x   ���9#��9l��9;��9A��9���9F��9���9���9F��9���9���9���9T��9N��9b��9���9��9���9��9���9���9���9(��9���93��9f��9��9���9���9x   x   !��9���9���9f��9���9>��9E��9���9���9���9���9P��9���9'��9���9:��9���9:��9���9��9���9���9���9��9���9���9��9���9���9���9x   x   ���9���9��9���9(��98��9{��9��9?��9j��9���9���9e��9���9���92��9���9v��9��9u��9.��9���9)��9���9���9��9���9���9o��9��9x   x   ���9;��9Z��9���9!��9���9@��9C��9���9���9&��9���9���9���9��9���9��9��9���9���9��9���9���9���9���9o��9���9���9��9���9x   x   ���9}��9���9	��9���9���9��9g��9��9Z��9���9��9��9���9���9i��9���9 ��9���9���9F��9r��9��9���9T��9���9K��9���9���9���9x   x   ��9��9��9���9���9/��9���9%��9���9���9l��9��9��9���9���9���9m��9��9N��9(��9���9���9���9���9���9���9w��9���9���9L��9x   x   ���9��9���9���99��9P��9���9b��9l��9���9��9E��9Y��9
��9���9N��9���9k��9���9B��9���9{��9E��9r��9���9��9+��9���9���9���9x   x   	��9���9���9���9���9P��9M��9*��9���9!��9��9���9���9��9r��9���94��9���9���9���9���9���9���9���9R��9���9���9���9��9r��9x   x   ���9���9=��9���9n��9���9(��9���9���9���9@��9���9��9���9���9���9��9+��9d��9���91��9���9���9��9(��9��97��9���9���9���9x   x   ���92��9T��9R��9���9S��9���9C��9���9L��9���9���9C��9/��9���9���91��9_��9��9���9q��9%��9}��9���9���9?��9 ��9��9���9���9x   x   ��9���9���9M��9$��9���9���9���9���9=��9���9v��9���9#��9p��9��9&��9���9���9���9G��9^��9���9���9��9���9B��9��9 ��9���9x   x   c��9#��9b��9,��9���9E��9���9y��9���9,��95��90��9P��9���9���9���9���9���94��9���91��9O��9~��9��9��9���9���9o��9!��9���9x   x   ��9���9p��9���9���9���9���9���9���9��9���9���9���98��9-��9���9&��9���9{��9���9p��9#��9v��9���9<��9���9���9[��9���9���9x   x   \��9���9���9��9���9N��9>��9,��9��9]��9a��9���9���9���9.��9���9���9���9G��9���9D��9��9	��9���9^��9���9���9v��9���9���9x   x   ���9k��9��9��9>��9���9���99��9���9d��9`��9x��9���9���9:��9���9���9���9���9��9���9���9���9L��9���9���9��9]��9���9���9x   x   
��9��9D��9���9���9���9x��96��9���9���9y��9���9���9���9��9h��9e��9w��9���9]��9���9��9_��9��9���96��9���9���9A��9���9x   x   ��9��9V��9���9��9A��9���9R��9���9���9���9���9C��9���9���9k��9���9p��9���9=��9]��9���9x��9���9���9���9��9��9���9���9x   x   ���9���9��9
��9���90��9$��9���96��9���9���9���9���99��9,��9���9/��91��92��9���9���9E��9���9~��9���9���9���9���9W��9���9x   x   ���9���9���9p��9���9���9s��9���9,��91��9=��9��9���9.��9���9���9���9m��9���9���9���9���9���9���9n��9���9���98��9���9���9x   x   h��9���9J��9���9���9���9��9���9���9���9���9i��9o��9���9��9r��9���9���9���9O��9���97��9���9���9��9V��95��9���9���9���9x   x   ���9m��9���93��9��9/��9#��9���9(��9���9���9h��9���90��9���9���9e��9?��9S��9���9���9t��9)��9@��9���9��9���9��9���9���9x   x   ��9��9k��9���9+��9c��9���9���9 ��9���9���9w��9s��9.��9q��9���9:��9c��9-��9���9'��9[��9_��9Z��9���9X��9��9���9���9 ��9x   x   ���9O��9���9���9`��9��9���92��9x��9G��9���9���9���9,��9���9���9V��9/��9L��9���9���9���9(��9���9���9���9���97��9��9���9x   x    ��9,��9D��9���9���9���9���9���9���9���9��9Z��9@��9���9���9M��9���9���9���9���9���9/��9{��9���9���9���9���9���9��9���9x   x   I��9���9���9���9.��9u��9G��92��9m��9B��9���9���9^��9��9���9���9���9*��9���9���9���9���9��9���9���9��9+��9F��9���9���9x   x   o��9{��9|��9���9���9'��9`��9P��9��9���9���9��9���9E��9��95��9r��9\��9���9/��9���9���9���9]��9���9���9���9���9���9���9x   x   ��9���9E��9��9���9|��9���9��9u��9��9���9]��9q��9���9���9���9&��9e��9,��9w��9��9���9 ��9���9���9���9;��9i��9���9��9x   x   ���9���9p��9���9��9���9���9��9���9���9O��9��9���9���9���9���9?��9\��9���9���9���9_��9���9���9���9���9���9���9���9?��9x   x   R��9���9���9T��9'��9���9��9��9<��9\��9���9���9���9���9p��9��9���9���9���9���9���9���9���9���9D��9F��9���9���9p��9���9x   x   ���9���9��9���9��9?��9���9���9���9���9���98��9���9���9���9S��9��9W��9���9���9��9���9���9���9G��9���9���9���9���9���9x   x   M��9x��9*��9���98��9��9E��9���9���9���9	��9���9��9���9���91��9���9��9���9���9)��9���9A��9���9���9���9���9���9���9���9x   x   ���9���9���9���9���9��9��9n��9_��9w��9Y��9���9��9���9=��9���9��9���97��9���9F��9���9i��9���9���9���9���9��9e��9B��9x   x   ���9���9���9��9���9���9 ��9 ��9���9���9���9>��9���9U��9���9���9���9���9��9��9���9���9���9��9p��9���9���9h��9K��9g��9x   x   ���9K��9���9q��9���9���9���9���9���9���9���9���9���9���9���9���9���9��9���9���9���9���9���9>��9���9���9���9F��9g��9=��9x   x   ͥ�9���9��9n��9���9<��9 ��9���9���9���9���9��9I��9��9ԫ�9���9��9۬�9ܫ�9w��9��9s��9��9���9���9Ш�9j��9ک�9��9ի�9x   x   ���9~��9z��9_��9���9���9Q��9��9ڭ�9���9d��9ج�9b��9���9���9i��9���9^��9}��9M��9���9b��9u��9@��9��9{��9d��9ƫ�9���9���9x   x   ��9~��93��9��9]��9���9W��9#��9:��9v��9	��9���9q��9M��9(��9���9#��9L��9��9���9 ��9���9���9���9V��9%��9r��9\��9O��9���9x   x   o��9_��9��9���9��9���9.��9��9��9���9^��9���9a��9���9ǭ�9���9��92��9���9N��9&��9Ѯ�9u��9i��95��9l��9s��9N��9���9���9x   x   ���9���9]��9	��9��9��9��9x��9��92��9��9��9���9���9���9��9��9y��9~��9��9ͫ�9��9���9���9���9���9��9ܬ�9��9ȭ�9x   x   ;��9|��9���9���9	��9��9H��9���9ڪ�9.��9ۤ�9u��9j��9/��9?��9���9l��9.��9I��9��9i��9��9���9���9ȫ�9G��9)��9\��9;��9ԩ�9x   x   ��9P��9[��90��9��9N��9(��9���9	��9���9��9٭�9.��9a��9���9���9j��9(��9I��9��9x��9���9y��9Ь�9��9p��9k��9)��9���9ƨ�9x   x   ���9��9&��9��9v��9���9���9���9S��9��9G��9B��9ʭ�9P��9ҭ�9���95��9@��9���9G��9���9��92��9Ħ�9G��9���9��9a��9­�9Ӫ�9x   x   ��9٭�95��9��9��9٪�9��9U��9p��9���9��9���9"��9���9��9=��9��9©�9��9n��9���9Z��9`��9���95��9}��9���9���9K��9���9x   x   ���9���9r��9���94��9/��9���9}��9���9���9���9��9���9��9ѭ�9��9���9G��9���9\��9��9r��9w��9=��9Ӭ�9٨�9x��9��9Ƭ�9���9x   x   ���9a��9��9d��9��9ڤ�9��9D��9��9���9���9���9ȫ�9&��9���9b��9#��9%��9:��9���9o��9���9+��9`��9g��9���9X��9��9���9Ϋ�9x   x   ��9֬�9���9���9��9s��9ڭ�9:��9���9x��9���9���9��9:��9��9]��9̮�9Ϊ�9���9̫�9s��9��9���9���9/��9>��9��9D��9��9��9x   x   L��9c��9p��9e��9���9j��90��9ɭ�9%��9���9ʫ�9%��9 ��9��9���9,��9_��9��9���9b��9��9��9A��9���9��9��9~��9���9��9U��9x   x   
��9���9N��9���9���9*��9c��9L��9���9��9#��9:��9��9���9���96��9g��9���9ܬ�9S��9��9��9 ��9/��9���9Ӭ�9:��9P��9z��9���9x   x   ӫ�9���9-��9˭�9���9?��9���9ϭ�9��9ѭ�9���9��9���9���9���9[��9Ԭ�9u��9���9X��9Ь�9r��9���9Ѭ�9ɩ�9��9n��9R��9V��9���9x   x   ���9n��9���9���9��9���9���9���9=��9��9g��9`��9&��98��9]��9���9���9L��9_��9���9U��9��9q��9��9F��9M��9���9n��9&��9��9x   x   ߫�9���9"��9��9��9k��9j��95��9��9���9 ��9ɮ�9\��9g��9Ӭ�9���9w��9��9���9��9���9���9���9خ�9���9q��9Ѭ�9��9���9��9x   x   ڬ�9[��9N��94��9|��91��9,��9D��9ĩ�9J��9!��9Ϊ�9 ��9���9y��9I��9��9���9���9Ȫ�9r��9��9���9Ϋ�9���9G��9��9>��9���9G��9x   x   ݫ�9z��9��9���9}��9D��9I��9���9��9���96��9���9���9ݬ�9���9_��9���9���9���9
��9��9'��9ɪ�9���9ŭ�9���9���9��9��9q��9x   x   v��9K��9���9P��9��9��9ޫ�9G��9r��9`��9���9ǫ�9a��9S��9Y��9���9��9̪�9��9Ϭ�9��9��9۪�9i��9D��9���9��9��9l��9y��9x   x   ��9���9 ��9$��9Ы�9j��9x��9���9���9��9t��9r��9��9��9Ь�9U��9���9p��9��9��9\��9A��9X��9��9���9L��9���9���9���9���9x   x   u��9e��9���9ή�9��9��9���9��9^��9p��9���9��9��9��9p��9���9���9~��9#��9��9?��9 ��9 ��9��9F��9���9Q��9ì�9���9���9x   x   ��9{��9���9x��9���9���9x��96��9g��9v��9)��9���9F��9 ��9���9q��9���9���9Ǫ�9ݪ�9V��9���9h��9���9>��9��9���9���9���9���9x   x   ���9?��9���9e��9���9���9ά�9¦�9���9>��9`��9���9���9,��9Ϭ�9��9خ�9˫�9���9g��9��9��9���9���9��9���9��98��93��9���9x   x   ���9	��9W��97��9���9ȫ�9��9K��97��9Ь�9c��90��9��9���9ȩ�9I��9«�9���9ȭ�9A��9���9H��9>��9��9��9��9
��9}��9��9ի�9x   x   Ө�9x��9(��9o��9���9I��9m��9���9~��9ݨ�9���9<��9��9Ҭ�9��9L��9q��9G��9���9���9J��9���9��9���9���9���9ة�9F��9?��9���9x   x   m��9b��9p��9n��9��9'��9j��9��9���9y��9T��9��9���9<��9q��9���9Ѭ�9��9���9��9���9R��9���9��9
��9ԩ�9��9���9���9���9x   x   ۩�9ǫ�9]��9N��9ެ�9[��9)��9a��9��9��9��9B��9���9P��9T��9n��9��9C��9��9��9���9Ŭ�9���9=��9~��9D��9���9���9m��9'��9x   x   ��9���9M��9���9��99��9���9ĭ�9H��9ɬ�9���9��9��9w��9T��9(��9���9���9��9l��9���9���9ª�95��9��9A��9���9g��9��9 ��9x   x   ֫�9���9���9���9ȭ�9֩�9Ǩ�9Ӫ�9���9���9ͫ�9��9T��9���9���9��9��9C��9k��9{��9���9���9���9���9ѫ�9���9���9'��9#��99��9x   x   @��9��9>��9d��9���9B��9o��9���9*��95��9��9.��9~��9���9Տ�9"��9���9���9l��9��9d��9���9c��9��9o��9͏�9Ж�9��9���9��9x   x   ��9���9��9��94��9���9��9��9b��9E��9��99��9��9���9j��9ב�9;��9
��9W��9L��9I��9���92��9��9U��9h��9���9ތ�9���9��9x   x   B��9��9���9l��9O��9���9���9ϐ�9ʒ�9���9Q��9��9p��9+��9L��9C��9��9��9_��9��9���9��9���9G��9̓�9z��9ג�9���9Ő�9'��9x   x   ^��9��9k��9s��9���9���9͋�9���9���9��9֐�9U��9���9Ԓ�9]��9V��9ܑ�95��9���90��9���9Ջ�9���9���9͐�9���9���9&��9%��9a��9x   x   ���98��9O��9���9'��9���9���9���9l��9���9n��9ˏ�9���9 ��9���9A��9���9
��9��9'��9���9:��9��9��9>��9���9@��9-��9���9���9x   x   C��9���9���9���9���9��9t��9��9��9ّ�9���9���9#��9��9$��9}��9H��9,��9ْ�9ɏ�9���9��9��9��9>��9��9���9���9���9i��9x   x   n��9��9���9ʋ�9���9v��9f��9{��9���99��9{��9Y��9ˑ�9���9���9���9e��9/��9���9a��9t��98��9��9N��9���9E��9L��9͋�9 ��9���9x   x   ���9��9͐�9���9���9��9~��9���9��9S��9̑�9y��9b��9���9j��94��9���9���9d��9ǐ�9���9���9���9��9.��9���9M��9���9���9��9x   x   (��9c��9˒�9���9n��9���9���9��9��9���9���9^��9ڐ�9`��94��9(��9p��9#��9���9��9I��9���9��9��9̑�9_��9#��9E��9���9 ��9x   x   4��9J��9���9��9���9ڑ�95��9R��9���9V��9v��95��9 ��9���9���9��9��9���9��93��9i��9v��9��9���9r��9ߒ�9���9}��9���9��9x   x   ��9"��9S��9Ԑ�9k��9���9|��9ˑ�9���9v��9���9o��9��9��9[��9��9���9���9���9���9���9V��9���9$��9���9ь�9e��9u��9܏�9c��9x   x   *��99��9��9T��9ȏ�9���9Y��9z��9d��9:��9q��9��9���9���9/��9ߐ�9���9X��9��9���9D��9���9���9��9&��9���9��9���9	��9Z��9x   x   ~��9��9m��9���9���9%��9ʑ�9b��9ِ�9 ��9��9���9��9B��9���9��9��9���9T��9��9���9O��9���9@��9&��9Ñ�9��9��9��9��9x   x   ���9Ɣ�9*��9В�9!��9��9���9 ��9a��9���9��9���9E��9��9���9s��9p��9f��9͐�9��97��9n��9c��9x��9C��9ԑ�9ג�9���9���9͐�9x   x   ׏�9e��9H��9\��9���9'��9���9m��96��9���9Z��9,��9���9���9֑�9ԑ�9��9i��93��9���9v��9œ�9���9r��9���9W��9��9;��9���9��9x   x   %��9ӑ�9A��9Q��9A��9}��9���95��9*��9	��9��9��9��9t��9ԑ�9���9���9{��9���9b��9���9x��9x��9ב�9<��9��9o��91��9���9Ȕ�9x   x   ���9@��9��9ܑ�9���9H��9c��9���9m��9��9���9���9��9q��9��9���9ĕ�9ד�94��9œ�9ϒ�9Z��9��9 ��9��9J��9q��9J��9x��9��9x   x   ���9��9��94��9��9'��9-��9���9��9���9���9]��9���9e��9j��9���9ߓ�9J��9<��9n��9O��9���9K��9���9Z��9^��9���9���9���9)��9x   x   n��9Z��9d��9���9��9ے�9���9m��9���9���9���9��9X��9̐�9-��9���92��98��9 ��9��9���9���9��9N��9��9���95��9��9Ƒ�91��9x   x   ��9M��9��9-��9+��9ȏ�9_��9ʐ�9��92��9���9Î�9��9��9���9c��9Ǔ�9n��9��9L��9���9���9���9��9{��9ϓ�9��9ԑ�9��9 ��9x   x   a��9H��9���9��9���9���9w��9���9F��9e��9���9B��9ޑ�94��9t��9��9Β�9L��9���9���9���9��9���9J��9���9��9
��9(��9r��9+��9x   x   ���9���9��9׋�9;��9��9>��9���9���9u��9U��9���9Q��9m��9Ǔ�9v��9X��9���9���9���9��9���9���9l��9-��9b��9���9R��9���9c��9x   x   `��9,��9���9���9��9��9��9���9���9���9���9���9���9c��9���9w��9��9L��9��9���9���9���9?��9ڐ�9���9U��9O��9��96��9���9x   x   ��9��9K��9���9��9��9O��9��9��9���9&��9��9:��9u��9t��9֑�9��9���9L��9��9N��9n��9ِ�9���9���9n��9J��9Z��9Ր�91��9x   x   m��9U��9Γ�9ǐ�9=��9?��9���9/��9ˑ�9q��9���9'��9&��9D��9���9<��9��9\��9���9{��9���90��9���9���9��9��9��9A��9o��9P��9x   x   Ώ�9i��9x��9���9���9 ��9E��9���9[��9��9ӌ�9���9đ�9ӑ�9Z��9��9H��9Y��9���9ϓ�9��9c��9S��9t��9��9]��9���9
��9O��9���9x   x   і�9���9ْ�9���9>��9���9O��9Q��9��9��9e��9��9��9ْ�9��9q��9r��9���95��9��9��9���9L��9L��9��9���9t��9C��9���9N��9x   x   }��9���9���9)��93��9���9Ћ�9���9D��9~��9t��9���9��9���97��9-��9I��9���9��9Α�9$��9S��9��9Y��9A��9��9A��9��9���9]��9x   x   ���9���9Ð�9%��9���9��9��9���9���9���9ݏ�9��9��9���9���9���9v��9���9Α�9��9t��9���94��9Ӑ�9p��9M��9ޒ�9���9U��9��9x   x   "��9��9'��9a��9���9l��9Ñ�9��9"��9��9`��9X��9��9ϐ�9��9Ɣ�9��9,��92��9���9*��9a��9���92��9P��9���9T��9\��9��99��9x   x   "}�9�v�93{�9|z�9Rv�9�}�9Oy�9�z�9�|�9�x�9�w�9)|�9�{�9�z�9�x�9Bz�9Sz�9a{�9s{�9	}�9?w�9y�9�|�9�x�9�y�9~�9�v�9Nz�9|�9�v�9x   x   �v�9�w�9I|�9ew�9�x�9�z�9u�9�x�9z�9�{�9�y�9�z�9x�9�y�9�z�9�z�97x�9�x�9~z�9�y�9[{�9qy�9oz�9u�9�y�9/x�9�w�9�{�9aw�9w�9x   x   .{�9I|�9y�9Gv�9�{�9�x�9Iy�9�w�9${�9�x�9{�9�y�9�v�9?y�9/w�9_z�9�w�9�y�9�z�9-y�9|�9�v�9}x�9�y�9�|�9v�9�y�9�|�9'{�9�w�9x   x   z�9fw�9Fv�9gy�9Hv�90{�9�|�9X}�9 y�9Ry�9{y�97y�9�|�9Fx�9Dw�91|�9�w�9`z�9�y�9�w�9~�9G}�9={�9nu�9�y�9�u�9w�9�z�9�|�9}�9x   x   Tv�9�x�9�{�9Gv�9�x�9�x�9�x�9�x�9�w�9�y�9�x�9�x�9�z�9�|�9�z�9!z�9Wy�9.x�9ly�9}x�9=x�9Iy�9�x�9Kv�9&|�9y�9?v�9�s�99{�9Ss�9x   x   �}�9�z�9�x�93{�9�x�9�u�9fy�9 }�9'y�9�{�9c{�9�w�9�|�9o}�9Uv�9�z�9�|�9�x�9o|�9*z�9~u�9�w�9�{�9xx�9az�9�}�9�v�9�z�9�z�9�v�9x   x   Ny�9u�9Iy�9�|�9�x�9gy�9)z�9%v�9"v�99v�9�r�9Bw�9�x�9w�9Ct�9Ru�9�v�92v�9z�9?y�9
z�9}�9�x�9�u�9*y�9z�9�{�9��9|�9�y�9x   x   �z�9�x�9�w�9Y}�9�x�9}�9)v�9�z�9j}�9y�9~�9�{�9�{�9�}�9 y�9/}�9Pz�9�v�9�|�9x�9�|�9�w�9�x�9.z�9
w�9�x�9�z�9ez�9 y�9,w�9x   x   �|�9z�9#{�9!y�9�w�9'y�9 v�9l}�9�w�9�y�9�|�9�z�9�}�9�x�9�x�9�}�9�u�9�x�9My�9y�9�{�9�y�9�|�9Py�9Gy�9�v�9.v�9�v�9py�9�x�9x   x   �x�9�{�9�x�9Py�9�y�9�{�98v�9y�9�y�9Vt�9�v�9�u�9=u�9Bz�9ow�9�v�9�{�9�x�9_x�9#y�9R{�9�x�9�y�9�{�9�y�9�y�98z�94y�9|�9z�9x   x   �w�9�y�9{�9}y�9�x�9d{�9�r�9~�9�|�9�v�94|�9�v�9�{�9�~�9�s�9cz�9�y�9mz�9�{�9�x�9�w�9�w�9�{�9�v�9�y�9U|�9�y�9�v�9�{�9zw�9x   x   %|�9�z�9�y�9>y�9�x�9�w�9Aw�9�{�9�z�9�u�9�v�9Z{�9�{�9|v�93w�9{y�9x�9y�9�z�9 }�9z{�9�y�9�x�9�w�9cx�9�w�94x�9_x�9�y�9K|�9x   x   �{�9 x�9�v�9�|�9�z�9�|�9�x�9�{�9�}�9;u�9�{�9�{�9�x�9`}�9�z�9e|�9�x�99x�9�{�9�{�95y�97w�9a{�9�w�9�s�9[x�9!{�9tw�99x�9|�9x   x   �z�9�y�9Cy�9Hx�9�|�9l}�9w�9�}�9�x�9Ez�9�~�9{v�9`}�9�{�9x�9�x�9�x�9*{�9�x�9�w�9�x�9@w�9{z�9?y�94y�9z�9�w�9sy�9�w�9�x�9x   x   �x�9�z�97w�9Ew�9�z�9Sv�9Et�9"y�9�x�9mw�9�s�94w�9�z�9x�9�w�9�z�9�y�9�z�9�y�9�{�9'{�9;x�9�z�9F|�9{�9�x�9"z�9�|�9ly�9�z�9x   x   Az�9�z�9^z�94|�9z�9�z�9Qu�9+}�9�}�9�v�9cz�9yy�9b|�9�x�9�z�9Pz�9�x�9�w�9\w�9�z�9k{�9Uy�9qy�9�y�9%y�9�{�9�z�9�v�9�w�9z�9x   x   Vz�97x�9�w�9�w�9Yy�9�|�9�v�9Wz�9�u�9�{�9�y�9x�9�x�9�x�9�y�9�x�9�w�97w�9�y�9�x�9Uw�9�x�9�z�9Yx�9�v�9y�9by�9x�9v�9zx�9x   x   a{�9�x�9�y�9_z�9-x�9�x�95v�9�v�9�x�9�x�9jz�9�x�99x�9,{�9�z�9�w�94w�9�}�9�z�9-y�9z�9�z�9�z�9{�9�x�9�z�9f}�9�w�9�x�92z�9x   x   p{�9~z�9�z�9�y�9ly�9n|�9z�9�|�9Ky�9^x�9�{�9�z�9�{�9�x�9�y�9Ww�9�y�9�z�9Hx�9{�9�w�9�u�9�v�9{�9�x�9�{�9%y�9Wv�9By�9�x�9x   x   }�9�y�9,y�9�w�9{x�9*z�9<y�9x�9y�9#y�9�x�9}�9�{�9�w�9�{�9�z�9�x�9,y�9{�9�w�9�w�9~x�9�w�9E{�9�w�9sx�9�{�9|�9�x�9�{�9x   x   Bw�9]{�9|�9~�95x�9u�9z�9�|�9�{�9T{�9�w�9x{�93y�9�x�9({�9i{�9Vw�9z�9�w�9�w�9�z�9�w�9'w�9�z�9mx�9Nz�9�z�9�x�9jx�9�{�9x   x   y�9py�9�v�9K}�9Iy�9�w�9
}�9�w�9�y�9�x�9�w�9�y�96w�9Bw�9=x�9Uy�9�x�9�z�9�u�9~x�9�w�9lv�9hz�9�w�9�y�9y�9�w�9�w�9�y�9�w�9x   x   �|�9mz�9}x�9;{�9�x�9�{�9�x�9�x�9�|�9 z�9�{�9�x�9`{�9|z�9�z�9qy�9�z�9�z�9�v�9�w�9*w�9gz�9�{�9ay�9�z�9
z�9�z�9nx�9{�9
z�9x   x   �x�9u�9�y�9ou�9Pv�9vx�9�u�93z�9Sy�9�{�9�v�9�w�9�w�9Dy�9F|�9�y�9[x�9{�9{�9A{�9�z�9w�9cy�9�|�98y�9�x�9�w�9?w�9|�9?y�9x   x   �y�9�y�9�|�9�y�9&|�9\z�9'y�9w�9Gy�9�y�9�y�9ax�9�s�93y�9{�9#y�9�v�9�x�9�x�9 x�9jx�9�y�9�z�94y�9^s�9�w�9y�9*y�9�x�9Xx�9x   x   ~�9-x�9v�9�u�9y�9�}�9 z�9�x�9�v�9�y�9R|�9�w�9Xx�9z�9�x�9�{�9y�9�z�9�{�9tx�9Kz�9y�9	z�9�x�9�w�9}�9�y�9�w�91x�9�x�9x   x   �v�9�w�9�y�9w�9>v�9�v�9�{�9�z�9/v�98z�9�y�98x�9${�9�w�9!z�9�z�9gy�9i}�9$y�9�{�9�z�9�w�9�z�9x�9y�9�y�9Pu�9�z�9\}�9\v�9x   x   Nz�9�{�9�|�9�z�9}s�9�z�9��9cz�9�v�95y�9�v�9_x�9pw�9ty�9�|�9�v�9x�9�w�9Zv�9|�9�x�9�w�9px�9@w�9)y�9�w�9�z�9<~�9�z�9s�9x   x   |�9`w�9){�9�|�99{�9�z�9|�9y�9py�9|�9�{�9�y�97x�9�w�9ky�9�w�9v�9�x�9?y�9�x�9jx�9�y�9{�9|�9�x�90x�9`}�9�z�9�{�9�|�9x   x   �v�9w�9�w�9}�9Os�9�v�9�y�9-w�9�x�9z�9yw�9I|�9|�9�x�9�z�9z�9{x�9/z�9�x�9�{�9�{�9�w�9	z�9;y�9^x�9�x�9[v�9s�9�|�9�v�9x   x   �f�9�c�9�a�9�a�9�e�9&a�9�c�9�a�9Oa�9�b�9�d�9�`�9	^�9�b�9a`�9�`�9�a�9�c�9j]�9a�9d�91b�9�a�9w`�9�d�9�b�9e�9Ma�9�a�9�c�9x   x   �c�9�^�9a�9�c�9�`�9ob�9�c�9c�9�a�9Ld�9c�9a�93d�9�b�9wb�97a�9Ua�9e�9�`�9	c�9$e�9ea�9�c�9xc�9�`�9�`�9/d�9La�9_�9�b�9x   x   �a�9a�9 f�9rc�9�a�9�a�9�d�9�a�9_�9ca�9�^�9vc�9�`�9�`�9�e�9�b�9�`�9�c�9_�9�`�9h_�9a�9�d�9c�9�a�9c�9�e�9�`�9�b�9e�9x   x   �a�9�c�9wc�9`f�9�b�9�b�96c�9�^�9�d�9Re�9�b�9�c�9�b�9�c�9�b�90b�9=c�9%c�9�e�9�c�9�_�9�c�9Aa�9sb�99f�9�c�99d�9�`�9�_�9�_�9x   x   �e�9�`�9�a�9�b�9c�9�b�9a�9�a�9�`�9�a�9c�9b�9�`�98^�9�`�9�c�9c�9>`�9b�9�a�9�_�9�c�9kc�9(b�9�a�9�_�9Lf�9�d�9�d�9pd�9x   x   %a�9pb�9�a�9�b�9�b�9Ob�9-e�9�a�91c�9�b�9�`�9�e�9d^�9�_�9�d�9I_�9�d�94c�9�`�9�e�9�a�9�a�9�b�9�a�9}b�9a�9bb�9Fc�9�c�9�b�9x   x   �c�9�c�9�d�97c�9a�90e�9a�9c�9]g�9 c�9�d�9�e�9b�9[e�9!g�97b�9vf�9�c�91a�9�e�9ma�9�b�9�d�9pc�90d�9T`�9�^�9C]�9A^�9W`�9x   x   �a�9c�9�a�9�^�9�a�9�a�9c�9�_�9b_�91g�9_^�9�_�9�_�9�]�9&g�9�_�9�_�9�c�9�`�9�`�9�_�9�a�9ec�95a�9�b�9hd�9�a�9#b�9�d�91c�9x   x   Qa�9�a�9_�9�d�9�`�90c�9[g�9d_�97a�9�`�9j_�9Kd�9�`�9L_�9�a�9�_�9f�9�c�9`b�9kd�9�^�9�a�9�a�9l`�9�d�9}e�9�_�9ae�9)d�9`�9x   x   �b�9Kd�9ea�9Ue�9�a�9�b�9c�9/g�9�`�9g�9�e�9Ld�9�g�9�a�9e�9d�9Vc�9�`�9�d�9�a�9e�9jb�9)b�9�a�9$c�9^a�9a�9Nc�9>b�9�b�9x   x   �d�9c�9�^�9�b�9	c�9�`�9�d�9a^�9p_�9�e�9#^�9�e�9�]�9s_�9f�9�_�9{c�9Rc�9S_�9qb�9Xd�9�^�9ld�90b�9�c�9b�9Xd�9�a�9�c�9a^�9x   x   �`�9a�9tc�9�c�9b�9�e�9�e�9�_�9Nd�9Nd�9�e�9�e�9�_�9�d�9e�9ub�9c�9�b�9a�9�`�9�a�9�c�9ub�9c�9uc�9�b�9�b�9�c�9Ld�9Sa�9x   x   
^�95d�9�`�9�b�9�`�9h^�9b�9�_�9�`�9�g�9�]�9�_�9Db�9{_�9�a�9�a�9na�9d�9;^�9�_�9�c�9id�9\b�9�c�9�c�9�d�9b�9.c�9�c�9�_�9x   x   �b�9�b�9�`�9�c�98^�9�_�9Ze�9�]�9N_�9�a�9n_�9�d�9{_�9x\�9�c�9xa�99b�9c�9�b�9�a�9�b�9#c�9c�9�d�9:d�9{b�9d�9Wc�9�a�9�b�9x   x   c`�9wb�9�e�9�b�9�`�9�d�9g�9#g�9�a�9	e�9f�9e�9�a�9�c�9�e�9�a�9a�9|c�9�b�9Ua�9�c�9Z`�9�_�9 a�9&`�9w`�94c�9�`�9�b�90d�9x   x   �`�98a�9�b�92b�9}c�9L_�98b�9�_�9�_�9d�9�_�9xb�9�a�9|a�9�a�9�`�9b�9�d�9�b�9�`�9�b�9�c�9b�9sb�9�c�9Pb�9}a�9�c�9�c�9�b�9x   x   �a�9Ra�9�`�9>c�9c�9�d�9qf�9�_�9f�9Oc�9xc�9�c�9pa�95b�9a�9b�9Td�9d�99c�9^a�9c�9Ic�9�c�9(b�9�c�9�a�9�a�9e�9cd�9�a�9x   x   �c�9e�9�c�9*c�9@`�95c�9�c�9�c�9�c�9�`�9Xc�9�b�9d�9c�9zc�9�d�9	d�9aa�9*a�9<d�9pb�9�a�9�b�9	c�9�c�9�a�9a�9�c�9e�9�b�9x   x   j]�9�`�9_�9�e�9b�9�`�91a�9�`�9`b�9�d�9U_�9a�9;^�9�b�9�b�9�b�9<c�9+a�9�^�9�c�9 d�9Dd�9�b�9�c�9�^�99b�9�b�9|b�9�c�9�b�9x   x   a�9c�9�`�9�c�9�a�9�e�9�e�9�`�9qd�9�a�9rb�9�`�9�_�9�a�9Pa�9�`�9]a�9;d�9�c�9{b�9�c�9$d�9�c�9Ve�9Cb�9�`�9"b�9@`�9�a�9{`�9x   x   d�9 e�9c_�9�_�9�_�9�a�9ma�9�_�9�^�9e�9Sd�9�a�9�c�9�b�9�c�9�b�9c�9pb�9d�9�c�9e�9�c�9�a�9xc�95e�9sa�9�c�9lc�9	c�9Pa�9x   x   1b�9fa�9a�9�c�9�c�9�a�9�b�9�a�9�a�9hb�9�^�9�c�9jd�9#c�9Z`�9�c�9Hc�9�a�9Dd�9'd�9�c�9Df�9Gb�9/a�9�c�9a�9Sc�9\d�9d�9�^�9x   x   �a�9�c�9�d�9Ba�9lc�9�b�9�d�9ec�9�a�9(b�9md�9wb�9]b�9c�9�_�9b�9�c�9�b�9�b�9�c�9�a�9Hb�9e�9�b�9�_�9nb�9�a�9
c�9�c�9:b�9x   x   v`�9xc�9c�9nb�9(b�9�a�9oc�94a�9k`�9�a�93b�9c�9�c�9�d�9a�9rb�9'b�9c�9�c�9We�9vc�9/a�9�b�9�`�9�d�9�d�9�b�9�a�9 b�93`�9x   x   �d�9�`�9b�97f�9�a�9b�9.d�9�b�9�d�9!c�9�c�9uc�9�c�9;d�9'`�9�c�9�c�9�c�9�^�9Bb�96e�9�c�9�_�9�d�9,c�9�b�9�c�9|c�9�c�9�c�9x   x   �b�9�`�9c�9�c�9�_�9a�9U`�9jd�9e�9\a�9b�9�b�9�d�9|b�9u`�9Ub�9�a�9�a�97b�9�`�9va�9a�9rb�9�d�9�b�9�b�9�`�9�e�9cd�9�^�9x   x   e�90d�9�e�9:d�9Mf�9`b�9�^�9�a�9�_�9 a�9Xd�9�b�9b�9d�92c�9za�9�a�9a�9�b�9 b�9�c�9Qc�9�a�9�b�9�c�9�`�9�_�9�a�9`�9b�9x   x   Pa�9Oa�9�`�9�`�9�d�9Dc�9D]�9$b�9_e�9Lc�9�a�9�c�9/c�9Zc�9�`�9�c�9	e�9�c�9zb�9B`�9pc�9Zd�9
c�9�a�9zc�9�e�9�a�9�[�9�c�9xe�9x   x   �a�9_�9�b�9�_�9�d�9�c�9C^�9�d�9)d�9Bb�9�c�9Ld�9�c�9�a�9�b�9�c�9`d�9e�9�c�9�a�9
c�9d�9�c�9%b�9�c�9cd�9`�9�c�9�c�9`�9x   x   �c�9�b�9	e�9�_�9pd�9�b�9Y`�91c�9`�9�b�9_^�9Ua�9�_�9�b�9/d�9�b�9�a�9�b�9�b�9x`�9Oa�9�^�9<b�93`�9�c�9�^�9b�9we�9`�9e�9x   x   �E�9GK�9xN�9^K�9�M�9XH�9
L�9�L�9�J�9�L�95M�9�L�9�N�9�J�9M�9�O�9�N�9�J�9�M�9�L�9�L�9�L�9PL�9�K�9M�9�I�9�K�9�J�9�M�9;K�9x   x   DK�9AR�91K�9�K�9�N�9�M�9EM�9�L�9M�9�H�9�L�95O�9DM�9�N�9M�9YK�9�M�9�M�9�O�9$M�9I�9xL�9$L�9nM�9�K�9VO�9mL�9�K�9�R�9J�9x   x   xN�9/K�9�I�9�K�9�J�9vM�9�I�9�O�9�N�9�L�9%M�9�L�9�M�9L�9-K�9�M�9�M�9+L�9�L�9L�9�N�9�O�9J�9WN�9�J�9�K�9�H�9�J�9�O�9VL�9x   x   ^K�9�K�9�K�9�I�9UN�94I�9KI�9M�9rM�9hL�9�J�9�K�9L�9�L�9oL�96K�93L�97K�9/M�9�L�9UM�9�I�9�G�9)O�9!I�9�L�9�L�9*J�9wJ�9�J�9x   x   �M�9�N�9�J�9ZN�9�M�9:M�9�N�98N�9�L�9~L�9�M�9�J�9DM�9�R�98M�9�K�9aM�97K�9tM�9�N�9�M�9PN�9�M�9	N�97K�9-M�9�M�9[N�9I�9�M�9x   x   ZH�9�M�9wM�98I�9:M�9]N�9gJ�9�K�9�J�9�H�9L�9�L�9L�9�L�9qL�9�J�9�J�9�J�9K�9�J�9�M�9lM�9'I�9vM�9�M�9�H�9�N�9�I�9�J�9�N�9x   x   	L�9FM�9�I�9II�9�N�9dJ�9
J�9�N�9�M�9K�9 L�9�M�9NN�9�L�9AM�9�J�9qL�9�O�9�I�9K�9_N�9�H�9�I�9�L�9�L�9GN�9�P�9M�9�O�9�N�9x   x   �L�9�L�9�O�9M�99N�9�K�9�N�9ML�9>K�9N�9J�9�N�9O�9BJ�9�M�9tK�9�L�91O�9*K�9N�9�M�9�O�9�L�9HL�9SN�9�I�9&N�9�N�9vI�9{N�9x   x   �J�9M�9�N�9pM�9�L�9�J�9�M�9BK�9M�9qN�9�K�9AK�9�K�9�M�9kM�9�K�9hL�9[K�97M�9#M�9$N�9�L�9�K�9�N�9J�9HK�9�P�9�K�9oI�9�N�9x   x   �L�9�H�9�L�9cL�9}L�9�H�9	K�9N�9qN�9�M�9�J�9J�9�N�9YO�9/L�9�K�9�I�9�K�9�L�9�L�9�I�9�L�9�N�9�I�9mJ�9�N�9]M�9�J�9�J�9ZO�9x   x   2M�9�L�9%M�9�J�9�M�9!L�9 L�9J�9�K�9�J�9cK�9lJ�9�I�9$K�9@M�9,K�9�M�9�J�9�L�9�L�9�L�9sO�9K�9�N�9BK�9I�9�L�9�M�9�I�9�O�9x   x   �L�94O�9�L�9 L�9�J�9�L�9�M�9�N�9<K�9J�9hJ�9�L�9�N�9{L�9SL�9�K�9GL�93L�9�O�9�L�9YM�9�J�9=K�9N�9�L�9L�9)M�9EM�9fK�96L�9x   x   �N�9CM�9N�9!L�9@M�9L�9RN�9O�9�K�9�N�9�I�9�N�9tN�9M�9�M�9�J�96N�9MM�9lN�9^N�9~K�9xL�9�I�9`J�9=N�9PK�9sI�9�J�9@L�9�N�9x   x   �J�9�N�9L�9M�9�R�9�L�9�L�9CJ�9�M�9TO�9#K�9|L�9M�9Q�9^M�9M�93N�9hJ�9�O�9]O�9�J�9�M�9�L�9zJ�9J�9�L�9vN�9|K�9O�9�N�9x   x   M�9M�9+K�9oL�99M�9pL�9=M�9�M�9jM�92L�9=M�9OL�9�M�9[M�9sJ�9EL�9$N�9 I�9NJ�9KL�9�K�9�M�9�M�9YL�9gM�9�M�9�K�9�J�9�K�9�I�9x   x   �O�9[K�9�M�93K�9�K�9 K�9�J�9yK�9�K�9�K�9.K�9�K�9�J�9M�9JL�9�O�9�M�9|K�9N�9�L�9�K�9�M�9wL�94M�9gN�9�J�9�M�9�N�9}I�9(N�9x   x   �N�9�M�9�M�92L�9aM�9�J�9rL�9�L�9eL�9�I�9�M�9DL�93N�91N�9'N�9�M�9�J�9�K�9@N�9\M�9�K�9}L�9�J�9K�9�L�9%M�9M�9xL�9iK�9~M�9x   x   �J�9�M�9'L�95K�9;K�9�J�9�O�93O�9]K�9�K�9�J�90L�9LM�9iJ�9I�9K�9�K�9MG�9�N�9SN�9J�9�J�9�K�9WJ�9CN�9=O�9G�9�K�9�J�9eH�9x   x   �M�9�O�9�L�9'M�9qM�9K�9�I�9)K�94M�9�L�9�L�9�O�9kN�9�O�9IJ�9N�9;N�9�N�9�M�96J�9\M�9�M�9�L�9�I�9{M�9�O�9�M�9N�9+L�9?O�9x   x   �L�9&M�9L�9�L�9�N�9�J�9K�9N�9!M�9�L�9�L�9�L�9_N�9ZO�9KL�9�L�9[M�9UN�95J�9�K�9iK�9K�9�L�9KK�9�L�9AM�9�M�9�J�9VN�9zO�9x   x   �L�9I�9�N�9WM�9�M�9�M�9aN�9�M�9#N�9�I�9�L�9YM�9|K�9�J�9�K�9�K�9�K�9J�9[M�9jK�9�F�9/K�9K�9+K�9M�9{J�9�K�9BL�9�K�9�L�9x   x   �L�9}L�9�O�9�I�9PN�9jM�9�H�9�O�9�L�9�L�9vO�9�J�9vL�9�M�9�M�9�M�9yL�9�J�9�M�9K�9-K�9oO�9K�9�J�9N�9tN�9XM�9`K�9�J�9?P�9x   x   LL�9&L�9J�9�G�9�M�9'I�9�I�9�L�9�K�9�N�9K�9;K�9�I�9�L�9�M�9uL�9�J�9�K�9�L�9�L�9K�9K�9�K�9)M�9|M�9�L�9"J�9QL�9�J�9yN�9x   x   �K�9jM�9XN�9*O�9N�9tM�9�L�9FL�9�N�9�I�9�N�9N�9^J�9{J�9[L�93M�9
K�9YJ�9�I�9MK�9-K�9�J�9'M�9�K�9�J�9�J�9zM�9�M�9|J�9�N�9x   x   M�9�K�9�J�9"I�97K�9�M�9�L�9VN�9J�9nJ�9CK�9�L�9?N�9J�9hM�9fN�9�L�9AN�9xM�9�L�9M�9	N�9yM�9�J�9�M�9�L�9�K�9K�9�I�9�N�9x   x   �I�9UO�9�K�9�L�9*M�9�H�9CN�9�I�9BK�9�N�9I�9L�9QK�9�L�9�M�9�J�9&M�9>O�9�O�9CM�9zJ�9uN�9�L�9�J�9�L�9�H�9�M�9�J�9J�97M�9x   x   �K�9jL�9�H�9�L�9�M�9�N�9�P�9&N�9�P�9`M�9�L�9%M�9oI�9sN�9�K�9�M�9M�9G�9�M�9�M�9�K�9WM�9 J�9zM�9�K�9�M�9�Q�9QN�9�P�9\N�9x   x   �J�9�K�9�J�9)J�9\N�9�I�9M�9�N�9�K�9�J�9�M�9EM�9�J�9~K�9�J�9�N�9xL�9�K�9N�9�J�9@L�9aK�9VL�9�M�9K�9�J�9PN�95L�9{J�9�O�9x   x   �M�9�R�9�O�9vJ�9I�9�J�9�O�9tI�9nI�9�J�9�I�9fK�9=L�9O�9�K�9~I�9gK�9�J�9/L�9UN�9�K�9�J�9�J�9{J�9�I�9J�9�P�9wJ�9	G�9�J�9x   x   ;K�9	J�9XL�9�J�9�M�9�N�9�N�9yN�9�N�9XO�9�O�99L�9�N�9�N�9�I�9(N�9zM�9cH�9BO�9yO�9�L�9AP�9vN�9�N�9�N�9<M�9_N�9�O�9�J�9�L�9x   x   B�9!8�9>6�9�9�94�9@9�96�9	8�98�9;7�9�6�9�7�9V:�9�8�9d8�9�3�9:�9�7�9P9�9�6�9�6�9�7�9%9�9�7�9o6�9�:�9J2�9q9�9X5�98�9x   x   "8�9�4�9�:�9�6�97;�9j9�96�98�9�8�9�8�9�7�9b5�9�3�9�6�9U8�9�6�9�6�94�9�6�9%8�9=8�9G8�9Q7�97�98�9z;�9�7�9[;�9:5�9{7�9x   x   ?6�9�:�9�9�9W9�9g6�9�9�9�8�9�6�9E9�9::�9�;�9\7�9�7�9[8�959�99�98�9Y6�9U:�9I:�9:�97�9�8�9�9�9�6�9�9�98�9�9�9�6�97�9x   x   �9�9�6�9S9�99�9�7�9<�9�;�9�7�93�9�4�9�7�9�7�9�:�9Y4�9�4�9�9�9}8�9�8�9�5�9A3�9�6�9�;�9~;�9u8�9�7�9�9�9�8�99�9�<�9�<�9x   x   4�99;�9d6�9�7�9�4�9�7�98�9�7�9�9�9�;�9�9�98�978�9�7�98�9f8�9�8�9^;�99�98�9�7�98�9z4�9�7�9{7�9n9�9h3�9h7�9<�9�6�9x   x   =9�9i9�9�9�9<�9�7�9R4�9�7�9:�9(8�9�9�9�<�9'6�978�908�9�6�9]<�9@:�9.8�9?:�9@8�9�3�9J8�9<�9-9�9i9�9�:�994�9�7�9�8�9&4�9x   x   6�96�9�8�9�;�98�9�7�9=�95�9�6�9�8�9�5�9e5�9�5�9�4�9�4�9i9�9�5�9�5�9�;�98�9�7�9G;�9)9�9�5�9E6�9A9�9P9�9x;�9�8�9�:�9x   x   8�98�9�6�9�7�9�7�9:�9!5�9�6�9�<�9�4�9<�9�7�9�8�9F=�9g4�9�<�9�6�95�9�:�9�7�9�7�9w6�9W8�98�96�96�9L5�9�5�9d5�9<6�9x   x   8�9�8�9B9�9|3�9�9�9$8�9�6�9�<�9�5�9w7�9�=�9�7�9�;�9o7�96�9�=�9�5�9�8�9w8�9b3�9�9�9B8�9�7�9�8�9<�9�7�9 3�9�8�9];�9_8�9x   x   =7�9�8�98:�9�4�9�;�9�9�9�8�9�4�9r7�9�1�98�99�9d2�9�7�9�3�9�8�9t:�97;�9\6�9�9�9�8�9�7�9p6�9�9�9�9�9,9�97�9�9�9�:�9k6�9x   x   �6�9�7�9�;�9�7�9�9�9~<�9~5�9<�9�=�98�9	B�9�7�9k<�9�<�9!6�9�;�9(9�9.8�9�:�9�7�96�9%8�9#7�94:�9�5�9�<�9[7�99�96�9�8�9x   x   �7�9a5�9_7�9�7�98�9(6�9e5�9�7�9�7�99�9�7�9�8�9k8�9�4�996�9 9�918�9�6�9�6�9�7�9E9�9�8�98�9�7�98�9�7�9�6�9P:�9�8�9>8�9x   x   Y:�9�3�9�7�9�:�958�998�9�5�9�8�9�;�9i2�9j<�9d8�9�5�9�8�9�7�9�9�98�9%4�9�8�9�5�97�9 ;�9�9�9�8�9�7�9�8�9�9�9�9�9�7�96�9x   x   �8�9�6�9Z8�9X4�9�7�9.8�9�4�9L=�9r7�9�7�9�<�9�4�9�8�97�9�4�9=9�9P6�9g8�9�6�97�9\7�9C7�9_9�9�7�9)8�9�9�9]7�9j8�9�6�9�4�9x   x   b8�9X8�939�9�4�98�9�6�9�4�9k4�96�9�3�9"6�996�9�7�9�4�9e8�9�7�9E9�9�:�9N7�9^;�9�8�9�6�9\9�9�;�9�8�9A6�9�8�9�9�9�9�9A;�9x   x   �3�9�6�9 9�9�9�9f8�9[<�9d9�9�<�9}=�9�8�9�;�99�9�9�9>9�9�7�944�9�7�9�:�9�5�9�8�9�9�9U5�9�6�9V7�9l6�9Z9�9�9�9�5�9�8�9c8�9x   x   :�9�6�98�9�8�9�8�9>:�9�5�9�6�9�5�9w:�9(9�958�98�9S6�9C9�9�7�96�9�9�9^7�9n6�9�7�9�:�9>:�9V9�9�7�9�5�9�7�9�9�9�6�9�7�9x   x   �7�94�9Z6�9�8�9`;�9(8�9�5�95�9�8�96;�9+8�9�6�9$4�9g8�9�:�9�:�9�9�9�;�907�9�5�9�:�9
:�93;�9�:�9�6�9�6�9�;�9W:�9M9�9�:�9x   x   P9�9�6�9X:�9�5�99�9D:�9�;�9�:�9x8�9^6�9�:�9�6�9�8�9�6�9M7�9�5�9a7�937�9F8�9:�9+9�9�4�9p8�9�9�9i8�9�7�9}6�96�9%9�9�6�9x   x   �6�9!8�9K:�9A3�98�9B8�98�9�7�9e3�9�9�9�7�9�7�9�5�9#7�9a;�9�8�9m6�9�5�9:�9�8�9o9�9;9�9�9�9�9�9�5�9�6�9N9�9::�9H5�9b6�9x   x   �6�9:8�9:�9�6�9�7�9�3�9�7�9�7�9�9�9�8�96�9C9�97�9^7�9�8�9�9�9�7�9�:�9+9�9n9�9F>�989�9:8�9S;�9�7�9
9�9�8�9_9�9$8�9c8�9x   x   �7�9D8�97�9�;�98�9J8�9C;�9w6�9<8�9�7�9#8�9�8�9 ;�9?7�9�6�9T5�9�:�9	:�9�4�9<9�9;9�9 5�9�:�9�9�96�9?7�96�9;9�9y8�9�8�9x   x   $9�9S7�9�8�9y;�9{4�9<�9)9�9X8�9�7�9p6�9 7�9�8�9�9�9a9�9Z9�9�6�9;:�9-;�9q8�9�9�9:8�9�:�9�9�9]7�98�9�9�9G;�9�9�97�9V5�9x   x   �7�97�9�9�9u8�9�7�9.9�9�5�98�9�8�9�9�92:�9�7�9�8�9�7�9�;�9[7�9V9�9�:�99�9�9�9T;�9�9�9`7�9�;�9|8�9o7�97�99�9�:�9�8�9x   x   n6�98�9�6�9�7�9z7�9f9�9D6�96�9<�9:�9�5�9
8�9�7�9$8�9�8�9k6�9�7�9�6�9i8�9�5�9�7�96�9!8�9}8�9�7�9�8�9�6�9U:�9�;�9�5�9x   x   �:�9z;�9�9�9�9�9n9�9�:�9@9�96�9�7�9+9�9�<�9�7�9�8�9�9�9B6�9V9�9�5�9�6�9�7�9�6�99�9B7�9�9�9k7�9�8�9d;�9S8�9$7�9�6�9n9�9x   x   O2�9�7�98�9�8�9k3�9=4�9N9�9L5�93�97�9[7�9�6�9�9�9^7�9�8�9�9�9�7�9�;�9|6�9P9�9�8�9#6�9I;�9�6�9�6�9T8�9�3�9$5�9D8�9a4�9x   x   o9�9\;�9�9�99�9f7�9�7�9v;�9�5�9�8�9�9�99�9T:�9�9�9i8�9�9�9�5�9�9�9W:�96�9::�9^9�999�9�9�99�9O:�97�9$5�9<�9�8�98�9x   x   Z5�995�9�6�9�<�9<�9�8�9�8�9e5�9`;�9�:�96�9�8�9�7�9�6�9�9�9�8�9�6�9L9�9$9�9F5�9%8�9u8�97�9�:�9�;�9�6�9F8�9�8�9:�9(=�9x   x   8�9x7�97�9�<�9�6�9)4�9�:�9;6�9`8�9m6�9�8�9;8�96�9�4�9A;�9f8�9�7�9�:�9�6�9b6�9b8�9�8�9W5�9�8�9�5�9m9�9`4�9 8�9%=�9�7�9x   x   ^ �9(&�9-#�9y&�9!)�9�&�9�$�9)(�9�%�9&�9.&�9�&�92'�9k'�9$�9\%�9�$�9g%�9�&�9�%�9F'�9'�9�%�93(�9�$�9}'�9(�9I&�9�"�9&�9x   x   (&�9x#�9�$�9(#�9+#�9$�9=&�9�&�9$�9�&�9�#�9*"�9b(�9%�9�&�9�%�9M&�9)�9z#�9�#�9%�9$�9 &�9�'�9e#�9�"�9.$�9v%�9�#�9?&�9x   x   +#�9�$�9�$�9�#�9�"�9�#�9�$�9�!�9"#�9}$�9I$�9�(�9�%�9#�9�)�9w"�9w%�9^'�9�#�9&%�9�#�9�"�9�#�9�"�9�#�9W$�93#�9E$�9/#�9'�9x   x   u&�9*#�9�#�9�*�9�$�9+$�9�#�9&�9�(�9U$�9,%�9<$�9�%�9�&�9S(�98%�9~%�9�%�9�#�9;)�9�$�9+$�9�$�9/%�9T)�9E$�94%�9|&�9!�9�9x   x   )�9+#�9�"�9�$�94$�9c%�9G#�9Q%�9"&�9u#�9� �9M#�9!&�9(!�9S%�9
#�9��9B$�99%�9�%�9�#�9�$�9�#�9%�9�#�9�!�9q'�9�&�90!�9�%�9x   x   �&�9$�9�#�9+$�9d%�9�(�9O&�9T �9c%�9�!�9�#�9H&�9&�9�%�9�'�9$�9�!�9�%�9p �9�&�9z(�9�%�9n$�9�"�9�#�9�(�9�&�9�%�9�&�9@&�9x   x   �$�9<&�9�$�9�#�9G#�9Q&�9d$�9�&�9�'�9�$�9�(�9](�9t)�9�'�9�&�9&�9u&�9z'�9�#�9&�9�#�9�#�9�$�9&�9�$�9�$�9B!�9\!�9-!�9$&�9x   x   ((�9�&�9�!�9&�9O%�9R �9�&�9�#�9�"�9�$�9�#�9��9� �9�$�9�$�9w"�9�$�9�&�9l!�9M%�9�%�9j!�9;'�9�(�9|$�9(�9�'�9a'�9&'�9�$�9x   x   �%�9$�9%#�9�(�9&�9^%�9�'�9�"�9�&�9�%�9V$�9#�9�"�9�&�9W&�9�"�9�&�9s%�9-%�9�(�9$�9�#�9�$�9r!�9�$�9�(�9�&�9�*�9$�9]!�9x   x   &�9�&�9~$�9V$�9w#�9�!�9�$�9�$�9�%�9&�9�$�9]&�9�%�9�%�91%�9�$�9�"�9#�9�%�9�#�9%&�9X'�9>%�9#�9�!�9$�9"�9�!�9�#�9�$�9x   x   0&�9�#�9E$�9&%�9� �9�#�9�(�9�#�9X$�9�$�9��9�$�9�$�9�#�9e(�9^#�9 �9]%�9�#�9�$�9�%�9#�9�&�9�$�9�#�9�'�9)%�9$�9�&�9$�9x   x   �&�9*"�9�(�9:$�9P#�9J&�9[(�9��9#�9[&�9�$�9#�9��9%(�9�&�9�#�9%�9�'�9�"�9'�9�%�9�$�9="�9T%�9�#�9�#�9�$�9#�9�$�9�$�9x   x   1'�9e(�9�%�9�%�9!&�9
&�9r)�9� �9�"�9�%�9�$�9��9�)�9�%�9�%�9�$�9q%�9R)�9�%�9�$�9P&�94%�9�#�9�'�9&�9'�9Y$�9T$�9�&�9�$�9x   x   m'�9%�9#�9�&�9%!�9�%�9�'�9�$�9�&�9�%�9�#�9&(�9�%�9�!�9�'�9�#�9�$�9'�9�#�9�&�9]$�9I$�9�#�9�#�95$�9$�9�#�9%�96&�9�!�9x   x   $�9�&�9�)�9S(�9U%�9�'�9�&�9�$�9_&�9/%�9f(�9�&�9�%�9�'�9�(�9J&�9$�9�#�9K%�9n%�9�#�9�%�9S$�9�#�9�#�99%�9m$�9*$�9R'�9�#�9x   x   `%�9�%�9z"�96%�9	#�9 $�9&�9s"�9�"�9�$�9^#�9�#�9�$�9�#�9G&�9�%�9�$�9c'�9�"�9�#�9p&�9�%�9$�9$�9y&�9Y&�9�#�9b"�9v&�9*%�9x   x   �$�9O&�9u%�9~%�9��9�!�9{&�9�$�9�&�9�"�9 �9%�9k%�9�$�9$�9�$�9,$�9$�9(%�9�&�9q&�9($�9$�9o#�9&�9{&�9�%�9�#�93%�9�$�9x   x   j%�9)�9\'�9�%�9A$�9�%�9y'�9�&�9r%�9#�9^%�9�'�9M)�9'�9�#�9e'�9$�9_%�9w$�90%�9�"�9�!�9�"�9#�9�%�9�#�9�%�9�$�9&�9$�9x   x   �&�9#�9�#�9�#�99%�9r �9�#�9o!�9/%�9�%�9�#�9�"�9�%�9�#�9O%�9�"�9(%�9w$�9�%�9�$�9L%�9_&�9x$�9:$�9�%�9>$�9�$�9�"�9z&�91$�9x   x   �%�9�#�9&%�97)�9�%�9�&�9 &�9K%�9�(�9�#�9�$�9'�9�$�9&�9j%�9�#�9�&�9/%�9�$�9�!�9s$�9D$�9�"�9�#�9�%�9�'�9�#�9%�98$�9%�9x   x   I'�9%�9�#�9�$�9�#�9y(�9�#�9�%�9$�9)&�9�%�9�%�9R&�9Y$�9�#�9p&�9m&�9�"�9M%�9p$�91"�9O$�9�$�9#�9^%�9J&�9�#�9N&�9�'�9�$�9x   x   '�9$�9�"�9,$�9�$�9�%�9�#�9m!�9�#�9['�9#�9�$�92%�9N$�9�%�9�%�9+$�9�!�9c&�9B$�9Q$�9&�9�"�9]$�9B&�9j&�9�"�9~#�9�$�9�"�9x   x   �%�9&�9�#�9�$�9�#�9q$�9�$�9:'�9�$�9@%�9�&�9;"�9�#�9�#�9S$�9$�9$�9�"�9{$�9�"�9�$�9�"�9�"�9i$�9�"�9�$�9�%�9�"�9�'�9�#�9x   x   3(�9�'�9�"�9.%�9%�9�"�9&�9�(�9r!�9#�9�$�9R%�9�'�9�#�9�#�9$�9r#�9#�9<$�9�#�9#�9^$�9j$�9E$�9F$�9�%�9�$�9A#�9�#�9"�9x   x   �$�9j#�9�#�9R)�9�#�9�#�9�$�9y$�9�$�9�!�9�#�9�#�9&�9:$�9�#�9z&�9&�9�%�9�%�9�%�9c%�9@&�9�"�9H$�9�&�9�$�9�%�9�!�9�#�9�#�9x   x   y'�9�"�9W$�9D$�9�!�9�(�9�$�9!(�9�(�9$�9�'�9�#�9'�9$�9<%�9\&�9z&�9�#�9>$�9�'�9N&�9e&�9�$�9�%�9�$�9]%�9�#�96)�9�(�9&�9x   x   (�90$�9.#�93%�9o'�9�&�9@!�9�'�9�&�9"�9.%�9�$�9V$�9�#�9k$�9�#�9�%�9�%�9�$�9�#�9�#�9�"�9�%�9�$�9�%�9�#�9�&�9H'�9q�95'�9x   x   F&�9x%�9F$�9~&�9�&�9�%�9[!�9d'�9�*�9�!�9$�9#�9T$�9%�9&$�9d"�9�#�9�$�9�"�9%�9O&�9}#�9�"�9@#�9�!�95)�9M'�9@#�9�%�9O&�9x   x   �"�9�#�9/#�9$�91!�9�&�9.!�9)'�9$�9�#�9�&�9�$�9�&�97&�9U'�9v&�90%�9 &�9{&�97$�9�'�9�$�9�'�9�#�9�#�9�(�9s�9�%�9(!�9i�9x   x   &�9?&�9'�9��9�%�99&�9"&�9�$�9\!�9�$�9$�9�$�9�$�9�!�9�#�9&%�9�$�9#$�94$�9%�9�$�9�"�9�#�9"�9�#�9	&�9/'�9K&�9g�9y'�9x   x   �	�9'�9��9>�9��9_�9<�9��9�9��9z�9f�9S�9`�9i�9��9��9�9��9��9��9��9M�9C�9��9E�9��93�9p�9�9x   x   #�9��9)�9q�9�9�9F�9��9!�9��9��9�9�9��9�9��9R�9��9��9�9��9��98�9�9r�9M�9�9��9��9?�9x   x   ��9+�9��9'�9��9-�9�9��9��9X�9�9��9��9��9w�9O�9t�9��9K�9��9��9��9{�9D�9��9��9��9��9��9F�9x   x   @�9q�9%�9��9�9-�9:�9��9/�9��9��9��9��9��9��9d�9��9Z�9'�9Z�9��9G�96�9��9��9b�9��9V�9;�9��9x   x   ��9�9��9�9 �9g�9+�9��9H�9��9��96�9�9��9��9��9��9(�9��96�9��9��9��9)�9^�9Q�9��9?�9��9��9x   x   a�9�9+�90�9c�9D�9]�9��9o�9�9��9��9��9��9�9��9��9�9W�9"�9��9��9c�9 �9�9��9�9]�9��9��9x   x   <�9E�9�99�9*�9]�9,�9��9Y�9{�9��9��9��9�9<�9��9��9��9��9�9k�9��9�9�9��9M�9��9��9!�9��9x   x   ��9��9��9��9��9��9��9��9��9j�9v�9��9��9��97�9��9$�9-�9�9��9��9��9*�9B�9q�9!�9��9Z�9h�9��9x   x   �9#�9��9.�9G�9q�9Y�9}�9��9(�9��94�9��9J�9��9z�9��9w�9��9#�9��9�9+�9��9��9 �9��9�9��9.�9x   x   ��9��9V�9��9��9�9{�9h�9*�9��90�9M�9��9��9��9��9\�9��9��9��9��9��9r�9��9��9`�9n�9��9��9��9x   x   x�9��9�9��9��9��9��9v�9��9/�9��9P�9d�9��9�9��9��9v�98�9��9��9��9�9�9��9�9��9*�9\�9Z�9x   x   i�9"�9��9��98�9��9��9��9-�9K�9M�9��9��9#�9y�9��9��9\�9X�9L�9O�9��9��9Z�9��9�9��9��9��9}�9x   x   P�9 �9��9��9�9��9��9�9��9 �9m�9��9��9��9��9w�9h�9��9��9[�9��99�9��9��9��9I�9?�9 �9l�9]�9x   x   a�9��9��9��9��9��9�9��9H�9��9��9"�9��9��9X�9_�9��9��9�9��9��9��9��9O�9K�9��9a�9T�9v�9�9x   x   h�9�9w�9��9��9�9;�96�9��9��9�9z�9��9X�9u�9�9��9\�9]�9c�9��9�9�9��9O�9��9��9��9��9��9x   x   ��9��9O�9e�9��9��9��9��9{�9�9��9��9y�9^�9�9��9��9��9��9U�9��9��9��9t�9��9X�9K�9@�9��9�9x   x   ��9R�9r�9��9��9��9��9�9��9]�9��9��9h�9��9��9��9y�9��9��9��98�90�9m�9��9��9Q�9��9��9��9��9x   x   �9��9��9]�9*�9 �9��92�9y�9��9t�9[�9��9��9X�9��9��90�99�9J�9��9u�9\�9j�9��9k�9��9��9y�9��9x   x   ��9��9J�9'�9��9W�9��9�9��9��96�9W�9��9�9\�9��9��97�9F�9��9I�9��9�9��9�9r�9�9�9��9	�9x   x   ��9!�9��9Y�98�9#�9�9��9#�9��9��9I�9Z�9��9d�9Y�9��9O�9��9��9��9 �9��9��9�9��9��9��9��9��9x   x   ��9��9��9��9��9��9m�9��9��9��9��9O�9��9��9��9��9;�9��9G�9��9��9��9��9��9��9�9��9��9i�9��9x   x   ��9��9��9D�9��9��9��9��9�9��9��9��99�9��9�9��90�9u�9��9�9��9��9\�9��9��9��9��9i�9��9��9x   x   L�9<�9{�99�9��9d�9�9,�9*�9o�9�9��9��9��9�9��9m�9]�9�9��9��9_�9�9�9��9��9��9��9��9��9x   x   D�9�9>�9��9&�9��9�9C�9��9��9�9]�9��9O�9��9q�9��9i�9��9��9��9��9�9��9b�9;�9�9��9��9��9x   x   ��9s�9��9��9^�9�9��9s�9��9��9��9��9��9H�9P�9��9��9��9�9�9��9��9��9`�9��9H�94�9��9i�9��9x   x   E�9L�9��9e�9Q�9��9M�9�9��9b�9�9�9J�9��9��9W�9S�9m�9s�9��9�9��9��98�9J�9��9E�9��9��9��9x   x   ��9	�9��9��9��9�9��9��9��9m�9��9��9C�9a�9��9J�9��9��9�9��9��9��9��9�91�9C�9n�9b�9I�9��9x   x   6�9��9��9V�9@�9_�9��9Y�9�9��9,�9��9�9Y�9��9B�9��9��9�9��9��9i�9��9��9��9��9a�9��9 �9V�9x   x   l�9��9��99�9��9��9!�9d�9��9��9\�9��9i�9t�9��9��9��9z�9��9��9g�9��9��9��9f�9��9H�9!�9��9^�9x   x   �9D�9E�9��9��9��9��9��9-�9��9Y�9|�9Y�9�9��9�9��9��9
�9��9��9��9��9��9��9��9��9V�9_�9��9x   x   ��9|�9���9��9��9H�9a�9��9��9q�9��9��9A�9��9N�9��9��9p�97�9��9��9f�9��9��9��9v�9�9��9���9{�9x   x   �9���9&�9��9��9��9$�9�9��9X�9� �9�9��9�9��9V�9��91�9�9� �9m�9*�9��9��9�9��9��91�9���92�9x   x   ���9$�9��9b�9��9��9X�9K �9�9��9��9�9�9��9��9��9��9/�9*�9��9<�9� �9�9��90�9b�9�9�9F��9���9x   x   ��9��9b�9l�9��9��9��9	��9���9��9���9� �9�9: �9b�9��9��9O��9��9 �9���9m�9��9�9�9G�9��9��9,�9i�9x   x   ��9��9��9��9�9q�9��9��9D�9��9��9w�9�9s�9� �9� �9c�9t�9
�9��9��9�9C�9��9`�9��9�9�9L�9�9x   x   K�9��9��9��9o�9X �9�9��9��9n�9R�9��9X�9@�9I�9��9�9��9+�9��9� �9��9c�9�9[�9��9��9���9���9�9x   x   b�9%�9U�9��9��9y�9�9z��9��9��9��9��9R��90�9��9I�9(�9R��9'�9��9��9��9��9��9�9��9�9��9>�9&�9x   x   ��9�9I �9
��9��9��9t��9
�9 �9� �9s�98�9L�9[�9�9)�9��9���9�9��9���9G �9��9��9|�9��9��9s�9��9L�9x   x   ��9��9�9���9D�9��9��9�9:��9d�9y �9/��9�9D�9h��9��9�9��9��9���9��9��94�96�9�9U�9��9�9R�9��9x   x   s�9X�9��9��9��9k�9��9� �9a�9��9� �9;�9�9�9U�9��9��9��9��9��9V�9J�9{��9��9��9��9�9��9� �9���9x   x   ��9� �9��9���9��9W�9��9q�9z �9� �9�	�9� �9'�9��9��9�9c�92��9>�9l�9~�9��9+��9��9+ �9n�9���9���9`��9��9x   x   ��9�9�9� �9x�9��9��9=�9+��9?�9� �9���9P�9,�9��9� �9�9��9��9R�9��9��9��9��9��9��9�9(�9��9��9x   x   C�9��9�9�9�9W�9N��9L�9� �9�9�9J�9N��9��97�9/�9��93�9��9:�9n�9��9��9�9��9q�9�9�9�9� �9x   x   ��9�9��97 �9|�9C�9+�9[�9B�9�9��9*�9��9��9j �9q	�9��9�9��9�9P�90�9`�9m�9��94�9�9��9;�9�9x   x   P�9��9��9[�9� �9K�9��9�9e��9V�9��9��97�9g �9��9�9��9~�9� �9t�9��9���9a�9(�9��9���9��9~�9���9��9x   x   	��9[�9��9��9� �9��9I�9.�9��9��9�9� �90�9p	�9�9���9�9��9X�9��9��9��9��9���9��9O�9�9"�9��9O�9x   x   ��9��9��9��9b�9�9&�9��9�9��9c�9�9��9��9��9�9��9�9 �97�9s�9��9&�9��9H�91�9���9�9�9��9x   x   n�95�91�9N��9s�9��9N��9���9��9��92��9��94�9��9~�9��9�9�9��9��9��9��98�9��9v�9Y�9��9��9:�9��9x   x   :�9�9)�9��9
�9'�9$�9��9��9��9;�9��9��9��9� �9W�9 �9��9��9T�9��9���9:�9r�9��9��9H �9��9t �9��9x   x   ��9� �9��9 �9��9��9��9��9���9��9n�9S�9:�9�9v�9��95�9��9O�9��9��9�9��9m�9_�9��9��9��9u�9�9x   x   ��9j�9:�9���9��9� �9��9���9��9Q�9~�9��9n�9O�9��9��9r�9��9��9��9f
�9��9��9�9��9��9��9{�9��9��9x   x   h�9*�9� �9k�9�9��9��9G �9��9I�9��9��9��9+�9���9��9��9��9���9�9��9���9o�9��9c�9���9� �9��9��9�9x   x   ��9��9�9��9B�9g�9��9��95�9}��9,��9��9��9`�9f�9��9%�96�9;�9��9��9n�9� �9G��9��9��9+�9�9���9���9x   x   ��9��9��9�9��9�9��9��96�9��9��9��9�9j�9&�9���9��9��9q�9o�9�9��9J��9��9�9��9��9���9r�98�9x   x   ��9�9/�9�9]�9\�9�9}�9�9��9+ �9��9��9��9��9��9I�9v�9}�9e�9��9a�9��9�9��9m�9S �9��9Q�9��9x   x   w�9��9a�9D�9��9��9��9��9V�9��9p�9��9q�95�9���9L�93�9[�9��9��9��9���9��9��9q�9U�9��9)�9��9�9x   x   �9��9�9��9�9��9�9��9��9�9���9�9�9�9��9}�9���9��9F �9��9��9� �9*�9��9S �9��9��9Z�9��9Q�9x   x   ��90�9�9��9�9���9��9s�9�9��9���9(�9	�9��9~�9$�9�9��9��9��9z�9��9�9���9��9+�9W�9��9���9� �9x   x   ���9���9J��9-�9J�9���9;�9��9R�9� �9a��9��9�9?�9���9��9 �9:�9s �9y�9��9��9���9s�9Q�9��9��9���9��93�9x   x   x�9-�9���9j�9�9�9'�9N�9��9���9��9��9� �9�9��9N�9��9��9��9 �9��9�9���9;�9��9�9Q�9� �93�9���9x   x   ���9���9���9i��9=��9<��9Z��9���9���9T��9���9��9i��9���9}��9m��9G��9���9
��9��9;��9K��9T��9a��9���9��9���9���9���9���9x   x   ���9���9���9���9���9��9���9R��9F��9���9���9 ��9���9���9���9���9��9���9���9=��9<��9Y��9E��9���9}��9���9���9l��9���9F��9x   x   ���9���9L��9%��9_��9Z��9���95��9���9���9���9���9f��9��9���9���9���9	��9���9���9���9n��9���9���9{��9���9���9��9���9���9x   x   i��9���9&��9&��9���9[��9e��9i��9?��9���9���9���9`��9���9l��9���9��9���9���9���9���9���9���9��9���9���9���9@��9��9���9x   x   :��9���9^��9���9v��9]��9B��95��9���9-��9���9���9���9���9T��9��91��9���9��9���9n��9s��9���9W��9H��9���9���9r��9���9��9x   x   7��9��9\��9\��9^��9/��9��9]��9��9���9[��9���9���9���9���9��9���9���9h��9H��9���9���9���9���9���9���9���9���9Q��9��9x   x   X��9���9���9g��9@��9��9���9U��9���9���9���9���9���9$��9d��9���9���9���9���9���9��90��9w��9p��9)��9���9���9M��9���9���9x   x   ���9Q��96��9h��94��9`��9R��9)��9%��9E��9V��9���9���91��9h��9-��9���9��9m��9a��9���9���9���9��9���9���9!��9v��9���9~��9x   x   ���9E��9���9@��9���9��9���9%��9v��9��9���9s��9���9S��9n��9���9���9@��9+��9(��9���9���9���9���9;��9M��9���9���9���9P��9x   x   S��9���9���9���9+��9���9���9D��9��9���9���9���9r��9���96��9���9/��9���9���9c��9a��9���9��9:��9���9"��9���9��9-��9���9x   x   ���9���9���9���9���9[��9���9W��9���9���9���9���9���9���9��9���9R��9v��9���9���9M��9D��9��9���9,��9p��9��9���9,��9���9x   x   ��9��9���9���9���9���9���9���9r��9���9���9���9���9w��9k��9���9���9���9���9Y��9���9���9���94��9a��9���95��9#��9!��9z��9x   x   k��9���9k��9f��9���9���9���9���9���9p��9���9���9��9���9z��9���9M��9@��9��9���9���9���9���9���9���9��9[��9g��9���9���9x   x   ���9���9��9���9���9���9$��93��9U��9���9���9{��9���9���9L��9���9G��9���9���9���9��9���9���9[��9���9���9���9���9���9���9x   x   y��9���9���9o��9P��9���9c��9g��9l��96��9��9k��9z��9L��9C��9��9-��9V��9���9���9���9���9���9���9.��9��9���9��9q��9��9x   x   j��9���9���9���9��9��9���9-��9���9���9���9���9���9���9��9���9L��9O��9w��9:��9Z��9���9���9���9-��9���9���9���9���9��9x   x   G��9��9���9��93��9���9���9���9���90��9S��9���9H��9H��90��9M��9{��9���9���9���9���9B��9B��9���9���9���9���9o��9���9���9x   x   ���9���9
��9���9���9���9���9��9B��9���9z��9���9?��9���9Y��9L��9���9c��9���9_��9e��9*��9���9E��9���9��9���9��9y��9���9x   x   ��9���9���9���9��9n��9���9o��9-��9���9���9���9��9���9���9t��9���9 ��9���9^��9��9���9n��9���9
��9G��9\��9 ��9���9���9x   x   ��9<��9���9���9���9H��9���9a��9%��9`��9���9Z��9���9���9���98��9���9b��9^��9a��9���9���9���9���9���9^��9��9l��9"��9���9x   x   ;��9>��9���9���9k��9���9	��9���9���9c��9K��9���9���9��9���9\��9���9h��9��9���9q��9���9��9���9���9j��9���9���9@��9���9x   x   J��9Y��9o��9���9x��9���93��9���9���9���9@��9���9���9���9���9���9A��9*��9���9���9���9'��9���9���9���9��9s��9W��9^��9n��9x   x   V��9A��9���9���9���9���9v��9���9���9��9��9���9���9���9���9���9D��9���9q��9���9��9���9��9���9���9o��9��9��9"��9P��9x   x   `��9���9���9��9W��9���9r��9��9���9=��9���93��9���9_��9���9���9���9E��9���9���9���9���9���9���9���9���9���94��9l��9���9x   x   ���9{��9|��9���9L��9���9*��9���9:��9���9.��9_��9���9���9(��9-��9���9���9
��9���9���9���9���9���9.��9���9f��9N��9`��9z��9x   x   ��9���9���9���9���9���9���9���9K��9!��9p��9���9��9���9��9���9���9��9E��9Y��9m��9��9m��9���9���9u��9p��9��9���9���9x   x   ���9���9���9���9���9���9���9 ��9���9���9!��93��9]��9���9���9���9���9���9]��9��9���9t��9��9���9j��9q��9���9Z��9���9���9x   x   ���9i��9��9=��9t��9���9Q��9x��9���9��9���9!��9l��9���9{��9���9p��9��9 ��9j��9���9Z��9��91��9N��9��9[��9���9���9���9x   x   ���9���9���9��9���9P��9���9���9���9,��9+��9"��9 ��9���9p��9���9���9{��9���9"��9>��9^��9%��9h��9_��9���9���9���95��9���9x   x   ���9G��9���9���9���9��9���9|��9O��9���9���9z��9���9���9��9��9���9���9���9���9 ��9q��9P��9���9w��9���9���9���9���9v��9x   x   s��9Y��9���9���9h��9��9o��9��96��9���9x��9	��9���9%��9���9���9P��9���9���9=��9U��9��9���9���9[��9���9>��9��9���9[��9x   x   V��9E��9_��9���9u��9���9@��9K��9W��9���96��9���9=��9'��9;��9���9���9���9���9���9j��9q��9���9��9a��9:��9���9���9���9o��9x   x   ���9`��9���9���93��9e��9���9���9[��9U��9���9���9#��9���9���9���9>��9m��9���9���9���9D��9���9���9���9}��9^��9���97��9��9x   x   ���9���9���9x��9N��9D��9���9���9��9��9V��9���97��9���9���9u��9q��9��9���9h��9���9e��9���9:��9���9��9��9���9���9���9x   x   h��9x��9/��9M��9'��9���9��9��9���9���9W��9Z��94��9���9���9���9
��9���9A��9���9���9 ��9���9!��9T��9���9���9���9 ��9���9x   x   ��9���9d��9E��9���9��9���9C��9���9���9��9��9���9a��9��9���9���9���9��9���9&��9���9���9���9��9��9���9���9���9���9x   x   o��9A��9���9���9��9���9h��9���9���9.��9���9A��9���9x��9���9��9���9Z��9[��9���9_��9��9K��9���9���9
��9���9a��9���9���9x   x   }��9I��9���9���9��9D��9���9x��9o��9���9C��9��9���9���9���9���9��9U��9���9��9_��9��9��9���9���9d��9���9���9���9���9x   x   9��9W��9]��9��9���9���9���9l��9���9���9���97��9���9���9��9���9p��9���9���9T��9��9���9���9���9���9���9G��9C��9���9*��9x   x   ���9���9P��9��9���9���9.��9���9���9��9<��9���9���9���9��9U��97��9���9���9���9N��9���9`��9���9%��9S��9H��9���9���9���9x   x   v��99��9���9X��9X��9��9��9D��9���9:��9&��9=��9���9���9{��9|��9���92��9x��9���9z��9s��9��9���9���9���9���9I��9s��9���9x   x   ��9���9���9���9Y��9��9C��9��98��9���9B��9���9���9b��9	��9(��9���9���9!��9���9y��9���9���9/��9���9Y��91��9���9F��9���9x   x   ���9:��9��96��95��9���9���9���9���9���9���9���9��9B��9]��9D��9%��9���9���9���9���9��9��9q��9���9��9��9��9~��9���9x   x   &��9*��9���9���9���9e��9z��9���9���9���9���9a��9@��9���9`��99��9[��9Z��9��9���9-��9���9���9��9��9���9���9��9���9���9x   x   ���9>��9���9���9���9��9���9���9��9��9x��9��9]��9^��9���9���9��9���92��9R��9���9���9���9"��9���9���9���9Q��9���9���9x   x   ���9���9���9w��9���9���9��9���9���9V��9y��9(��9H��97��9���9���9���9^��9���9���9���9���9A��9���97��9���9z��9*��9���9���9x   x   U��9���9:��9s��9��9���9���9��9n��96��9���9���9(��9Z��9��9���9���9{��9���9���9���9���90��9���9���9���9���9���9���9\��9x   x   ���9���9q��9��9���9���9[��9U��9���9���91��9���9���9Z��9���9`��9z��9��9��9���9���9���9<��9"��9���9���9!��9l��9��9���9x   x   ���9���9���9���9@��9��9Z��9���9���9���9x��9��9���9��92��9���9���9��9���9���9U��9��9���9��9���9���9���9��9���9��9x   x   >��9���9���9h��9���9���9���9��9S��9���9���9���9���9���9S��9���9���9���9���9���9���9z��9��9 ��9���9���9���9���9���9���9x   x   S��9k��9���9���9���9)��9e��9]��9��9L��9{��9x��9���9,��9���9���9���9���9U��9���9k��9���9@��9"��9���9���9l��9���9���90��9x   x   ��9o��9E��9c��9��9���9��9��9���9���9v��9���9
��9���9���9���9���9���9��9|��9���9���9���9T��9)��9+��9���9d��9h��9���9x   x   ���9���9���9���9���9���9N��9��9���9[��9��9���9���9���9���9F��9/��9<��9���9��9@��9���9���9���9y��9���9���9���9���9!��9x   x   ���9��9���9?��9'��9���9���9���9���9���9���92��9r��9��9&��9���9���9��9��9!��9"��9S��9���9i��9���9b��91��9p��9���9���9x   x   \��9_��9���9���9V��9��9���9���9���9#��9���9���9���9 ��9���9:��9���9���9���9���9���9*��9z��9���9���9[��9���9���9��9���9x   x   ���9>��9|��9��9���9~��9��9e��9���9S��9���9X��9��9���9���9���9���9���9���9���9���9/��9���9b��9S��9��9��9s��9S��9���9x   x   <��9���9^��9��9���9���9���9���9K��9J��9���95��9��9���9���9|��9���9��9���9���9o��9���9���95��9���9��9���9���9��9D��9x   x   ��9���9���9���9���9���9_��9���9B��9���9I��9���9��9��9S��9*��9���9j��9	��9���9���9f��9���9p��9���9o��9���9b��9���9V��9x   x   ���9���96��9���9���9���9���9���9���9���9q��9D��9���9���9���9���9���9��9���9���9���9f��9���9���9��9R��9��9���9���90��9x   x   \��9s��9���9���9���9���9���9���9+��9���9���9���9���9���9���9���9\��9���9��9���90��9���9"��9���9���9���9G��9V��94��9���9x   x   R��9C��9���9T��9���9f��9���9'��9���9���9��9���9��9���9���9���9���9���9���9+��9��9A��9��9Z��9m��9���9���9���9���9E��9x   x   F��9W��9���95��9-��9���9^��9���9���9���9���9>��9���9���9O��9J��9���9 ��9���9���9���9t��9r��9���9��9���9���9:��9|��9���9x   x   ���9���9n��9��9l��9@��9���9���9���9X��9q��9f��9H��9��9-��9<��9���9���9&��9���9���9%��9���9���9���9���9Z��9��9���9$��9x   x   V��90��9��9���9���9���9���96��9���9x��9���9���9,��9��9��9���9��9���9R��9��9!��9���9v��9���9(��9���9���9��9A��9r��9x   x   ���9,��9o��9���9���9��9G��9���9���9��9���9���9���97��90��9���9���9<��97��97��9 ��96��9���9���9���9j��9$��9
��9��9(��9x   x   g��9���9;��9���9��9R��9s��9��9F��9J��9G��9���9��9���9���9\��9]��9#��9��9h��9���9d��9��9���9���9L��9��9e��9���9���9x   x   ���9_��9���9���9J��9o��9���9~��9}��9���9���9���9 ��9���9
��9���9���9���9K��9���9c��9���9B��9d��9j��9���9��9���9���9���9x   x   '��9���9���98��9���9��9��9���9���9���9���9���9��9���9���9���9���9/��9���9���9���9���9��9���9S��9Y��9���9���9���9���9x   x   ���9���9���9���9���9I��9��9���9���9D��9���9��9?��9���9���9d��9���9���9��9S��9O��9��9���9���9G��9 ��9���9���9'��9���9x   x   ���9���9W��9z��9��9H��9���9���9D��9���9���9���9u��9U��9���9��9v��9���9��9���9���9���9���9��9��90��9���9���9���9E��9x   x   ��9���9m��9���9���9G��9���9���9���9���9���9���9��9���9���9u��9���9M��9&��9���9���96��9���9[��9��9N��9���9j��9���9j��9x   x   ���9A��9d��9���9���9���9���9���9��9���9���9���9X��9|��9���9���9���98��90��9��9d��9��9u��9���9C��9U��9���9��9y��9r��9x   x   ��9���9M��9-��9���9��9��9��9A��9q��9���9U��9P��9���9s��9���9/��9���9���9d��9���9��9y��9\��9I��9���9-��9��9���9<��9x   x   ���9���9��9��9:��9���9���9���9��9Y��9���9|��9���9���9���9��9g��9,��93��9���9F��9l��9���9��9���9���9|��9���9���9���9x   x   ���9O��9,��9��93��9���9��9���9���9���9���9���9u��9���9]��9���9Q��9���9���9>��9s��9j��9��9���9���9X��9���9���9%��99��9x   x   ���9M��99��9���9���9Y��9���9���9d��9 ��9s��9���9���9��9��9���9���9���9���9���9���9F��9���9���9���9%��9���9���9t��9���9x   x   ���9���9���9	��9���9`��9���9���9���9z��9���9���9.��9e��9T��9���9��9���9���9���91��9|��9`��9I��9���9���9���9O��9 ��9���9x   x   ���9 ��9���9���9?��9'��9���92��9���9���9K��96��9���9+��9���9���9���99��90��9���9���9���9���9���9��9���9���9���9���9 ��9x   x   ���9���9!��9U��98��9 ��9K��9���9��9��9$��90��9���94��9���9���9���90��9���9���9H��9B��9S��9���9v��9B��9��9���9���9���9x   x   *��9���9���9��98��9f��9���9���9T��9���9���9��9b��9���99��9���9���9���9���9���9��9���9���9!��9���9U��9���9���9T��9!��9x   x   ��9���9���9 ��9��9���9c��9���9Q��9���9���9`��9���9J��9u��9���9.��9���9H��9��9N��9N��9���9���9��9$��9���9���9���90��9x   x   A��9t��9(��9���95��9a��9���9���9��9���9:��9���9��9o��9o��9I��9{��9���9A��9���9M��9���9@��92��9'��9���9V��9��9p��9���9x   x   ��9p��9���9w��9���9��9E��9��9���9���9���9w��9x��9���9��9���9^��9���9P��9���9���9@��9���9N��9���9P��92��9���9l��9���9x   x   Z��9���9���9���9���9���9b��9���9���9��9Z��9���9Y��9��9���9���9I��9���9���9��9���94��9O��9���9���9���9���9���9���9���9x   x   l��9
��9���9(��9���9���9k��9S��9G��9��9��9E��9I��9���9 ��9���9���9��9p��9���9��9$��9���9���9[��9e��95��9t��9���9E��9x   x   ���9���9��9���9i��9P��9���9Z��9���9/��9P��9Y��9���9���9[��9!��9���9���9?��9X��9 ��9���9P��9���9c��9f��9��9���9���9f��9x   x   ���9z��9Y��9���9#��9	��9��9���9���9���9���9���9)��9���9���9���9���9���9	��9���9���9S��9.��9���94��9��9���9d��9���9���9x   x   ���99��9��9��9��9g��9���9���9���9���9i��9��9��9���9���9���9P��9���9���9���9���9��9���9~��9u��9���9e��9��9G��9���9x   x   ���9y��9���9B��9	��9���9���9���9'��9���9���9~��9���9���9#��9v��9 ��9���9���9U��9���9u��9n��9���9���9���9���9C��9���9���9x   x   G��9���9%��9v��9(��9���9���9���9���9F��9j��9p��99��9���9;��9���9���9���9���9&��91��9���9���9���9E��9h��9���9���9���9��9x   x   ���9���9@��9��9���9���9���9���9M��9���9K��9��9v��97��9���9r��9|��9-��93��9��9���9���9��9y��9@��9f��9���9T��9e��9���9x   x   ���9f��9���9���9���9���9W��9���9���9]��9���9���9��9��9;��9���9���9>��9���9w��9���9���9���9���9 ��9��9a��9���9��9���9x   x   @��9���9���9���9A��9;��9?��9N��9Y��9���9d��9���9���9���9��9C��9���9���9���9	��9���9L��9��9A��9��9��9��9���9m��9���9x   x   ��9���9��9���9x��9���9���9���9���9 ��9'��9Q��90��9)��9=��98��9���9���9t��9���9���9���9#��9r��9���92��9���9���9��9���9x   x   ���9���9?��9z��9[��9T��9���9��9���9���9���9T��9���9���9��9E��9"��9'��9O��9���9���9��9���9���9���9���9���9\��9���9@��9x   x   ���9���9:��9���9S��9���9S��9]��9���9��9���9���9���9��9���9���9W��9���98��9;��9w��9u��9J��9���95��9`��9���9]��9���9N��9x   x   ���9Z��9B��9���9���9R��9���9:��9<��9���9?��9���9��9���9���9���9@��9���9T��9���93��9���9-��9���9��9���9���9<��9y��9z��9x   x   ���9���9M��9���9��9`��98��9���9���9���9���9���9���9���9��9;��9��9���9���9��9���9���9���9l��9��9^��9 ��9���9=��9��9x   x   P��9���9W��9���9���9���96��9���9���9��9z��9%��95��9i��9"��9p��91��9���9���9S��9���9K��9,��9R��9���9���9���9f��9#��9N��9x   x   ���9[��9���9 ��9���9��9���9���9���91��9 ��9��9h��9u��9h��9���9o��9���9���9���9+��9���9���9���9���9���9���9P��9S��9���9x   x   J��9���9h��9*��9���9���9A��9���9v��9��9}��9��9e��9U��9���9<��9���9b��9r��9x��9O��9���9���9���9���9��9n��9���9D��9|��9x   x   ��9���9���9O��9Q��9���9���9���9��9��9��9���9���9���9��9���9#��9>��9���9���9f��9?��9���9���9���9X��9?��9���9���9���9x   x   y��9��9���9.��9���9���9��9���96��9g��9f��9���9T��9���9���9���9O��9���9���9��9���9���9I��95��9E��9|��9���9q��9
��9���9x   x   :��9��9���9%��9���9��9���9���9m��9y��9U��9���9���9U��9���9���9���9���9��9���9���9��9��9���9��9X��9���9,��9���9c��9x   x   ���98��9��9=��9��9���9���9��9��9c��9���9��9���9���9P��9'��9��9���9H��9E��9���9���9=��9.��9���9���9���9���9��99��9x   x   v��9���9G��98��9F��9���9���9>��9q��9���9;��9���9 ��9���9)��9���9���9���9M��9
��9���9��9L��9~��9��9x��9���9���9���9���9x   x   {��9���9���9���9$��9V��99��9 ��92��9n��9���9#��9P��9���9��9���9���9���9]��9|��9���9���9���9���9o��9���9*��9��9���9B��9x   x   /��99��9���9���9"��9���9���9���9���9���9d��9@��9���9���9���9���9���9X��9���9#��9���9$��9[��9/��9���9[��9���9���9~��9���9x   x   8��9���9���9t��9J��9<��9V��9���9���9���9t��9���9���9��9L��9N��9\��9���9���9���9���9/��9��9���9��9���9��9���9���9,��9x   x   ��9x��9	��9���9���9=��9���9��9P��9���9y��9���9��9���9G��9	��9}��9%��9���9��9���9���95��9[��9R��9���9���9���9��92��9x   x   ���9���9���9���9���9u��93��9���9���9,��9O��9i��9���9���9���9���9���9���9���9���9��9���9 ��9���9���9j��9J��9���9A��9���9x   x   ���9���9K��9���9��9z��9���9���9I��9���9���9=��9���9
��9���9��9���9"��9,��9���9���9���9���9���9���9���9��9H��9���9���9x   x   ��9���9��9!��9���9K��9*��9���9+��9���9���9���9J��9���99��9N��9���9\��9��95��9$��9���9���9	��9���9���9���9`��9C��9��9x   x   z��9���9C��9q��9���9���9���9k��9Q��9���9���9���97��9���9.��9���9���91��9���9^��9���9���9��9���9���9��92��9���9���9���9x   x   A��9���9��9���9���96��9��9��9���9���9���9��9G��9��9���9��9n��9���9��9Q��9���9���9���9���98��9���9���9���94��9���9x   x   e��9��9��9/��9���9\��9���9a��9���9���9 ��9R��9~��9U��9���9{��9���9]��9���9���9o��9���9 ��9��9���9C��9s��97��9���9|��9x   x   ��9d��9��9���9���9���9���9!��9���9���9q��9;��9���9���9���9���9&��9���9��9���9M��9��9���93��9���9m��9��9[��9���91��9x   x   T��9���9���9���9\��9`��9<��9���9e��9R��9���9���9r��9+��9���9���9��9���9���9���9���9N��9[��9���9���98��9\��9[��9���9���9x   x   e��9��9n��9��9���9���9w��9?��9"��9R��9B��9���9
��9���9��9���9���9���9���9��99��9���9H��9���94��9���9���9���9��9���9x   x   ���9���9���9���9A��9N��9z��9	��9N��9���9y��9���9���9d��96��9���9B��9���9,��97��9���9���9��9���9���9~��93��9���9���9���9x   x   ���9���9���94��9=��9���9���9���9��9M��9_��9���9o��9���9���9O��9j��9���9���9���9���9��9F��9 ��9��9���9���9��9i��9���9x   x   ���9���9��9���9)��9���9���9���9x��9<��9���9W��9���9���9���9���9���9���9��9���9���9���9��9���95��9���9���9���9���9���9x   x   ���9��9��9���9���9���9D��9���9��9���9>��9���9��9���9���9���9~��9���9X��9 ��92��9���9 ��9���9���9b��9p��9���9B��9B��9x   x   /��9���9���9���9���9���9 ��9��9G��9P��9��9J��9w��9D��9���9��9���9/��9���9y��9���9W��9o��9&��9��9���9���9���9|��9���9x   x   ;��9(��9���9���9��9p��9&��9���9D��9U��9���9���9���9���9@��9W��9��9���9��9���9���9���92��9���9���9)��9��9,��9{��9i��9x   x   ���9��9���9���9r��9���9���9���9���9��9���9���9��9���9��9���91��9n��9n��9���9���9��9���9���9S��9��9B��9���9n��98��9x   x   ���9���9B��9 ��9$��9���9<��9��9���9���9���9x��9Q��9���9���9M��9���9���9���9��9��9���9,��9���9���9��9n��9���9���9A��9x   x   ���9���9���9��9���9���9��9���9���9��9���9%��9��9���9���9z��9l��9	��9���9K��9R��9��9���9q��9}��9L��9���9���9��9&��9x   x   ��9|��9��9J��9B��9���9���9���9���9��9��9C��9���9/��9|��9���9q��9���9`��9���9���9W��9���9n��9?��9f��9���9i��9���9���9x   x   M��99��9���9N��9T��9��9���9��9��9���9j��9���9���9l��9��9���9'��9A��9���9]��9���9���9n��9H��9���9���9���9���9$��9���9x   x   a��9���9<��9��9���9���9���9���9��9l��9���9w��9���9���9��9���9��9���9J��9���9i��9/��9��9���9c��9���9���9���9��9���9x   x   ���9Y��9���9J��9���9���9s��9!��9G��9���9y��9���94��9W��9���9���9"��9���9��9���9s��9��9:��9.��9���9���9m��9_��9���9E��9x   x   m��9���9��9z��9���9��9I��9��9���9���9���97��9���9���9p��9���9D��9���9���9���9���94��9I��9c��9���9���9��9n��9���9��9x   x   ���9���9���9F��9���9���9���9���9-��9k��9���9[��9���9���9p��9���9��9U��9���9n��9��9���9���9 ��9���9@��9*��9!��9M��9���9x   x   ���9���9���9���9<��9��9���9���9|��9"��9��9���9m��9m��9���9���9���9���9���9F��9���9i��9���9U��9���9���9���9A��9L��9���9x   x   P��9���9���9��9[��9���9R��9~��9���9���9���9���9���9���9���9O��95��9���9>��9���9���9��9��9���9���9���9���9���9���9���9x   x   o��9���9z��9���9
��94��9���9n��9q��9&��9��9 ��9C��9��9���99��97��9H��9[��9w��9���9��9���9��9<��9���9%��9J��9���9���9x   x   ���9���9���9/��9���9q��9���9��9���9?��9���9���9���9W��9���9���9K��9M��92��9���9���9��9��9���9���9���9��9���9��9��9x   x   ���9���9U��9���9��9m��9���9���9d��9���9I��9��9���9���9���9?��9Z��91��9m��91��9,��9���9���9���9t��9)��9��9���9	��9���9x   x   ���9���9���9}��9���9���9��9I��9���9^��9���9���9���9j��9I��9���9w��9���9-��9��9��9#��9+��9���9k��9���9���9b��9y��9���9x   x   ���9���93��9���9���9���9��9S��9���9���9h��9v��9���9��9���9���9���9���90��9��9���9*��9���9���9���9���9)��9���9#��9\��9x   x   ��9���9���9W��9���9��9���9��9T��9���92��9��94��9���9l��9��9��9
��9���9&��9*��9���9���9/��9���94��9���9U��9���9���9x   x   H��9��9���9n��9.��9���9/��9���9���9s��9 ��97��9H��9���9���9��9���9��9���9'��9���9��9���9d��9���9��9���9���9 ��98��9x   x   ��9���9���9)��9���9}��9���9r��9m��9I��9���90��9c��9��9T��9~��9��9���9���9���9���9,��9a��9���9L��9h��9���9���9 ��9���9x   x   ��97��9���9��9���9Q��9���9{��9>��9���9_��9���9���9���9���9��9>��9���9t��9l��9���9���9���9L��9{��9���9*��9y��9C��9���9x   x   ���9���9]��9���9*��9��9��9L��9h��9���9���9���9���9A��9���9���9���9���9+��9���9���90��9���9i��9���9���9|��9���9���9��9x   x   ���9���9p��9���9��9D��9o��9���9���9���9���9m��9��9(��9���9���9&��9 ��9 ��9���9&��9���9���9���9-��9y��9a��9���9U��9���9x   x   ��9���9���9���9+��9���9���9���9i��9���9���9]��9j��9"��9C��9���9K��9���9���9b��9���9U��9 ��9���9z��9���9���9=��9S��9N��9x   x   h��9���9B��9���9y��9n��9���9��9���9"��9��9���9���9I��9J��9���9���9��9��9y��9#��9���9���9���9E��9���9U��9V��9��9H��9x   x   ���9���9>��9���9j��98��9B��9%��9���9���9��9J��9��9���9 ��9���9���9��9���9���9`��9���95��9���9���9 ��9���9N��9E��9��9x   x   ��98��9͹�9���9���9$��9���9���96��9Y��9/��9���9��9���9���9���9i��9d��9���9��9��9���9��9Z��9E��9y��9��9X��9��9]��9x   x   4��9���9i��9���9º�9$��9���9L��9��9��9���9��9A��9R��9���9C��9���9���9���9l��9���9��9ƻ�9���9H��9��9u��9��9���9Թ�9x   x   й�9m��9G��9$��9��93��9>��9���9B��9ʺ�9x��9߽�9��9��9&��99��9n��9b��9}��9ۻ�9z��9��9Ժ�9V��9g��9���9x��9���9��9q��9x   x   ���9���9"��9u��9���9^��9ɼ�9ٻ�9!��9��9׺�9��9���9��9��9���9���9��9���93��9T��9R��9|��9Ƚ�97��9��9w��9.��9��9ھ�9x   x   ���9º�9���9���9߸�9��9���9p��9}��9��9B��9��9v��9��9��9;��9Ž�9��9Ի�9���9Ժ�9���9˸�9?��9���9E��95��9��9���9-��9x   x   !��9!��92��9]��9��9ǻ�9���9��9���9��9x��9=��9r��9��9º�9���9���9u��9���9;��9���9��9���9���9ƻ�9���95��9��9g��9���9x   x   ���9���9?��9ȼ�9���9���9O��9��9x��9���9��9��9��9Z��9���9��9���9��9��9<��9'��9ؼ�9���9+��9���9���9��9���9���9���9x   x   ���9O��9���9ػ�9n��9޹�9��9ѿ�9���9���9(��9��9��9���9߹�9���9߿�9��9���9���9���9���9ۺ�9��9���9ɷ�9m��9��9��9E��9x   x   4��9��9@��9 ��9���9���9y��9���90��9���9��9x��9U��9Һ�9B��9ռ�9l��9A��9ֺ�9��9���9Ժ�9º�9%��9���9N��9��9���9���9]��9x   x   Y��9���9˺�9��9��9��9���9���9���9��9��9̻�9���9��9��9V��9��9R��9��9���9��9Q��9]��9��9��9��9^��9���9'��9���9x   x   /��9���9t��9Ժ�9@��9w��9��9(��9��9��9&��9��9���9��9Ҹ�9ȼ�9J��9ܻ�9P��9i��9G��9`��9���9���9$��9���99��94��9���9r��9x   x   ���9��9߽�9��9��9;��9��9��9{��9ǻ�9��9Ǹ�9��9���9@��9J��9t��9���9���9A��9b��9���9A��9��9���9��9��9%��9ܽ�9j��9x   x   ��9C��9��9���9s��9r��9��9��9X��9���9���9��9���9��9���9��9ϻ�9��9��9$��9���9��9 ��9��9��9��9ѽ�9ҹ�9,��9׼�9x   x   ���9P��9��9��9��9��9]��9���9Ժ�9��9��9���9��9��9\��91��9޺�9���9���9���9^��9f��9���9޹�9q��9���9���9��9_��9'��9x   x   ���9���9&��9��9��9���9���9��9@��9��9и�9@��9���9_��9a��9���9P��9��9���9���9��9���9��9ս�9x��9���9���9���9��9���9x   x   ���9D��9:��9���9<��9��9��9��9ϼ�9R��9ļ�9H��9��96��9���9W��9��9n��99��9&��9��9��9;��9<��9'��9���9P��9��9���9���9x   x   h��9���9n��9���9ƽ�9���9��9߿�9g��9��9M��9v��9ѻ�9��9R��9!��9+��9��9���9��9)��9b��9���9u��9���9,��9���9���9���9���9x   x   `��9���9d��9��9��9r��9��9��9@��9S��9ܻ�9���9��9���9��9l��9��9��9��9x��9d��9��9��9y��9���9���9y��9v��9k��9��9x   x   ���9���9y��9���9Ի�9���9��9���9Ӻ�9��9P��9���9��9���9���94��9���9 ��9R��9۹�96��9Y��94��9���9:��9��9ܼ�9)��9Ľ�9��9x   x   ���9o��9ڻ�92��9���9=��9?��9���9��9��9j��9E��9"��9���9���9'��9��9|��9۹�9U��9���9Y��9���9���9л�9���9���9ƾ�9��9Ȼ�9x   x   ��9���9z��9T��9պ�9���9(��9���9���9��9C��9^��9���9a��9��9��9'��9i��94��9���9R��9���9��9���9e��9P��9���9V��9D��9��9x   x   ���9��9��9R��9���9��9ؼ�9���9Ժ�9P��9`��9���9��9i��9���9߻�9b��9��9X��9V��9���9��9R��9w��9���9���9���9��9��9ݻ�9x   x   ��9Ż�9պ�9��9̸�9���9���9غ�9���9W��9���9B��9���9���9��98��9���9��91��9���9��9R��9��9r��9���9+��9l��9P��9��9ڻ�9x   x   [��9���9S��9ƽ�9:��9���9%��9��9)��9��9���9��9���9��9ս�97��9|��9}��9���9���9���9{��9t��9���9���9���9���90��9���96��9x   x   D��9I��9f��97��9���9̻�9���9���9���9!��9%��9���9��9r��9y��9#��9���9���98��9λ�9d��9���9���9���9��9 ��9���9ʿ�95��9��9x   x   v��9��9���9��9E��9���9���9ķ�9J��9��9���9��9��9���9���9���90��9���9��9���9O��9���9+��9���9!��9E��9/��9غ�9���9���9x   x   ��9s��9w��9w��90��95��9��9m��9��9_��97��9��9н�9���9���9N��9���9t��9޼�9���9���9���9l��9���9���94��9���9���9��9L��9x   x   X��9��9���9-��9��9��9���9��9���9���97��9(��9ӹ�9$��9¾�9��9���9x��9,��9ʾ�9X��9��9T��9-��9ɿ�9ܺ�9���90��9ٸ�9`��9x   x   ��9���9��9��9���9i��9���9��9���9%��9���9ݽ�9*��9]��9��9���9���9h��9ý�9���9E��9��9��9���92��9���9��9ܸ�9o��9d��9x   x   Y��9Թ�9o��9ܾ�9*��9���9���9A��9^��9���9p��9j��9Ѽ�9%��9���9���9���9��9��9û�9��9ۻ�9޻�92��9��9���9H��9^��9b��9���9x   x   ���9���9~��9��9��9���9)��9���9���9���9���9;��9d��9B��9)��9^��9���9{��9���9��9���9?��9���9���9`��9޵�9���9��9��9���9x   x   ���9���9��9D��9���9@��9m��9Ҵ�9T��9���9���9t��9?��9Բ�9���9[��9���9_��9��9R��9ͷ�9?��9{��9��9��9ӷ�9���9���9���9{��9x   x   |��9��9J��9g��9���9���9��9D��9���9-��9(��9O��9_��9b��9���9���9���9T��9��9���9��9t��9���9_��9]��9ó�9���9G��9���9��9x   x    ��9C��9f��9���9��9<��9F��9���9��9x��9���97��9J��9��9���9���9��9p��9c��9��9��9��9���9;��9u��9f��9"��9l��9��9f��9x   x   ��9���9���9��9|��9e��9��9 ��9p��9���9γ�9%��9���9���9��9��9˲�9N��9T��9q��9��9���9ϲ�95��9ɰ�9*��95��9}��9��9Ȱ�9x   x   ���9@��9���9;��9e��9���9ѵ�9 ��9R��9̱�9���9���9_��9���9��9��9߲�9���9���9}��9���9/��9���9��9H��9��9��9{��9i��9���9x   x   *��9n��9��9C��9���9е�9?��9���9F��9+��9Ƶ�9N��9\��99��9ߵ�9���9���9��9���9���9/��9���9	��9z��9j��92��9��9���9��9��9x   x   ���9Ӵ�9D��9���9��9#��9���9���96��9r��9^��9t��9D��9}��9��9��9���9���9���9���9ߴ�9���9e��9J��9ֵ�9���9���90��9̶�9��9x   x   ���9S��9���9	��9l��9R��9D��90��9���9)��9���9��9	��9[��9��9���9���9\��9y��9���9z��9g��9]��9���9.��9��9���9̶�9��9���9x   x   ���9���9.��9w��9���9˱�90��9t��9,��9���9ܵ�9��9���9V��9���9v��9ǳ�9���9!��9���9��9s��9j��91��9���9ڴ�9��96��9���9̳�9x   x   ���9���9,��9���9ҳ�9���9ŵ�9[��9���9ݵ�9i��9ߵ�9	��9���9O��9���9���9���9��9���9w��9˳�9��9o��9��9��9���9γ�9߶�9��9x   x   9��9v��9P��95��9(��9���9O��9p��9޶�9��9ߵ�9.��9��9ش�9>��9��9��9ѵ�9��9Z��9{��9Y��9���9ʰ�9��9��9K��9���9���9|��9x   x   d��9=��9a��9I��9���9[��9Z��9@��9��9���9	��9��9F��9��9\��9U��9]��9f��9��9x��9���9l��9B��9���9���9���9}��9״�9��9W��9x   x   F��9ղ�9e��9��9���9���97��9|��9X��9P��9���9ִ�9��9��98��9׵�9ղ�9���9���9I��9��9u��9ڸ�9��9̴�9���9C��9��9���9���9x   x   +��9���9���9���9��9��9��9��9��9���9Q��9B��9]��98��9��9ϱ�94��9w��9I��9H��9y��9?��9!��9���9ܴ�9���9+��9���9���9��9x   x   ]��9\��9���9���9��9��9���9��9���9x��9���9��9P��9ӵ�9α�9
��9���9b��9���9��9���96��9��9���9��95��9Դ�9W��9Q��9կ�9x   x   ���9���9���9��9̲�9��9���9���9���9ʳ�9���9��9[��9Ӳ�9/��9���9]��9��9���9#��9��9���9I��9��9 ��9ʷ�9���9���9i��9���9x   x   ~��9^��9T��9o��9L��9���9��9���9[��9���9���9ҵ�9e��9���9u��9b��9��9��9 ��9���9���9��9v��9@��9_��9n��9��97��9˳�9��9x   x   ���9��9��9c��9S��9���9���9���9z��9#��9��9��9��9 ��9M��9���9���9��9k��9P��9X��9��9���9i��9B��9��9���9-��9���9���9x   x   ��9P��9���9��9s��9y��9���9���9���9���9���9\��9v��9F��9H��9��9 ��9���9O��9���9���9���9��9��9Q��9��9��9���9C��9���9x   x   ���9̷�9��9��9��9���9-��9ߴ�9z��9��9y��9~��9���9��9y��9���9��9���9W��9���9���9}��9���9&��9,��9c��9���9÷�9з�9��9x   x   C��9A��9t��9��9���90��9���9���9h��9w��9γ�9W��9i��9r��9?��9;��9���9��9��9���9}��9&��9���9��9b��9���9���9��9"��9f��9x   x   ���9}��9���9���9ϲ�9¶�9	��9f��9`��9j��9��9���9D��9ٸ�9��9��9G��9p��9���9��9���9���9���9ִ�9��9*��9���9��9Ƿ�9��9x   x   ���9��9_��9>��94��9 ��9{��9N��9���9,��9n��9˰�9���9��9���9���9��9=��9i��9��9&��9��9ٴ�9c��9���9���9@��9���9P��9x��9x   x   c��9��9[��9w��9ư�9J��9k��9ص�9*��9���9��9��9���9˴�9ܴ�9��9���9\��9B��9O��9*��9]��9 ��9���9���9H��9���9���9!��9~��9x   x   ݵ�9ѷ�9���9d��9$��9ߵ�90��9���9��9ݴ�9��9��9���9���9���99��9˷�9q��9��9��9d��9���9&��9���9M��9ٸ�9��9ٶ�9:��9��9x   x   ���9���9���9$��99��9��9ݳ�9���9���9��9���9I��9���9@��9*��9մ�9���9��9���9��9���9���9���9>��9���9��9
��9Ų�92��9���9x   x   ��9���9I��9n��9��9|��9���91��9ȶ�96��9γ�9���9ִ�9��9���9V��9���96��9)��9���9���9��9��9���9���9ն�9ò�9��9{��9���9x   x   ��9���9���9��9��9k��9}��9ж�9��9���9߶�9���9��9���9���9U��9p��9ϳ�9���9I��9ӷ�9��9Ƿ�9S��9"��9:��91��9~��9R��9���9x   x   ���9}��9��9g��9ʰ�9���9��9��9���9ͳ�9��9z��9[��9���9��9ѯ�9���9|��9���9���9��9c��9��9y��9���9��9���9���9���9���9x   x   ��9���9���9���9&��9��94��9���9���9��9���9��9���9���9��9p��9���9A��9��9��9��9���9��9���9Ĭ�9���9.��9���9��9���9x   x   ���9���9���9���9���9߱�9q��9���9���9��9|��9ȭ�9ˬ�9���9���9���9���9C��9��9c��9M��9j��9��9]��9ڰ�9��9���9���9���9���9x   x   ���9���9��9@��9��9��9A��9��9{��9���9���9R��9D��9)��9���9N��9Ϯ�9$��91��9b��9��9���9���9���9_��9̮�9}��9^��9��9���9x   x   Ĳ�9���9?��9��9.��9��9L��9���9R��9]��9���9j��90��9��9I��9l��9���9��9���9��9���9��9���9X��9 ��9���9���9\��95��9��9x   x   #��9��9��9.��9_��9���9֮�9��9���9X��9��9��9ٮ�9ҭ�9L��9��9ձ�9Ӱ�9���9~��9Ю�9$��9��9e��9���9���9]��9K��9|��91��9x   x   ��9��9��9��9���9���9%��9]��92��9ū�9Ư�9���9��9ݯ�9	��9V��9���9"��9)��9ͮ�9���9E��9j��9��90��9��9���9��9>��9��9x   x   5��9p��9C��9L��9Ԯ�9"��9���9���9U��9���9��9G��9��9���9°�9p��9l��9d��9b��9[��9��9T��9���9��9��9���9=��9#��9���9ʰ�9x   x   ���9���9��9���9��9[��9���9���9��9��9k��9��9��9���9)��9s��9 ��9���9��9��9��96��9��9I��9Į�9&��9���9)��9֮�9L��9x   x   ���9���9{��9T��9���92��9W��9���9���9˰�9]��9��9���9Ӱ�9���9���9���9���9���9��9���9׮�9���9��9��9_��9��9���9t��9���9x   x   ��9��9���9]��9W��9ƫ�9���9��9˰�9���9G��9E��9V��9���9���9��9
��9���9خ�91��9��9��9��9Y��9*��9���9T��9h��9;��9ΰ�9x   x   ���9y��9���9���9��9���9��9j��9_��9K��9ޭ�9>��9���9��9���9���9@��9��9?��9��9D��9ͮ�9I��9��9_��9��9%��9���9���9T��9x   x   ��9ɭ�9Q��9i��9��9��9H��9��9��9I��9;��9+��9v��9~��9¯�9���9���9���9��9���9��9���93��98��98��9��9Į�9���9��9׭�9x   x   ���9Ȭ�9G��9-��9خ�9��9��9��9���9V��9���9v��9߮�9N��9Я�9���93��9���9��9���9���9���9���9��9]��9ʰ�9���9���9���9���9x   x   ���9���9*��9��9ҭ�9ݯ�9���9���9ְ�9���9
��9��9N��9ˬ�9P��9ܰ�9��9@��9��9̰�9+��9@��9���9���9ʮ�9��9#��9��9��9j��9x   x   ��9���9���9G��9N��9��9���9'��9���9���9���9¯�9ϯ�9Q��9���9Q��9Ӯ�9���9h��9í�9���9���9���9*��9Ǫ�9��9���9G��9��9���9x   x   p��9���9S��9l��9��9U��9n��9j��9���9��9���9���9���9ް�9T��9���92��9t��9-��9���9ر�9K��9D��9I��9���9/��9d��9��9���9M��9x   x   ���9���9Ү�9 ��9Ա�9���9m��9���9���9��9@��9���94��9��9׮�95��9���9X��9���9v��9���9Ǯ�9���9Э�9���9���9��9:��9���9���9x   x   D��9D��9 ��9߯�9Ӱ�9 ��9c��9���9���9���9��9���9���9C��9���9t��9W��9k��9>��9+��9!��9���9'��9���92��9��9c��9o��9=��9w��9x   x   ��9��9/��9���9���9*��9c��9��9���9ۮ�9?��9��9��9��9h��9,��9���9@��9m��9e��9S��9���9��9)��9���9m��9=��9��9g��9h��9x   x   ��9_��9c��9��9{��9ʮ�9[��9��9��92��9��9���9���9ǰ�9���9��9y��9-��9g��9���9��9���95��9���9���9/��9��9���9���9k��9x   x   ��9L��9��9���9Ү�9���9!��9��9��9��9B��9��9���9-��9���9ձ�9���9!��9T��9��9���9Ʈ�9��9	��9Ū�9İ�9_��9-��9���9���9x   x   ���9h��9���9��9&��9G��9T��98��9Ү�9��9ɮ�9���9���9B��9���9H��9ɮ�9���9���9���9Ȯ�9^��9
��9���9Ƭ�9_��9���9A��9c��9	��9x   x   ���9��9���9���9��9f��9���9��9|��9��9L��94��9���9���9���9A��9���9(��9��91��9��9
��9T��9`��9a��98��9���9��9��9ٯ�9x   x   ���9Y��9���9Y��9f��9��9��9G��9|��9`��9��97��9��9���9*��9G��9ͭ�9���9+��9���9��9���9a��9|��9į�9I��9���9���9���9J��9x   x   Ĭ�9ذ�9_��9!��9���9,��9��9���9��9+��9^��9;��9[��9Ǯ�9ɪ�9���9���92��9���9���9ʪ�9Ǭ�9c��9ʯ�9]��9լ�9^��9��9���9]��9x   x   ���9��9ˮ�9���9���9��9���9*��9\��9���9��9��9ɰ�9��9��9.��9���9��9i��9)��9Ű�9\��98��9G��9Ӭ�9���9��9��9��9#��9x   x   ,��9���9��9���9^��9���9<��9���9��9R��9%��9î�9���9(��9��9e��9��9g��9?��9���9_��9���9���9���9^��9��9N��9ݰ�9S��9U��9x   x   ���9���9`��9Y��9G��9��9"��9+��9���9h��9 ��9���9���9��9F��9��97��9l��9��9���9+��9@��9��9���9��9��9��9���97��9��9x   x   ��9���9��97��9{��9?��9���9خ�9r��9=��9���9
��9���9۱�9��9���9���9=��9c��9���9���9h��9|��9���9���9��9R��96��9߭�9A��9x   x   ���9���9���9��9.��9��9ɰ�9J��9���9а�9W��9ӭ�9���9h��9���9P��9���9w��9i��9i��9���9��9ׯ�9J��9]��9!��9U��9��9?��9��9x   x   "��9&��9���9ҩ�9c��9ۨ�9T��9��9��9D��9���9��9��9y��9/��9Ө�9���9���9���9��9Q��9���9ݧ�9���9Ĭ�9���9��9*��9���9��9x   x   #��9Ϭ�9W��9���9h��9���9��9_��9o��9r��9Ȭ�9��9s��9��9\��9���9��9k��9���9Z��9���9��9���9���9��9)��9N��9��9���9���9x   x   ���9U��9~��9���9���9���9:��9a��9'��9��9x��9��9"��9̦�9`��9���9���9��9f��9���9���9(��9:��9ب�9���9���9���9���9_��9Э�9x   x   ҩ�9���9���9ͬ�9b��9��9:��9Ȫ�9ī�9X��9צ�9F��9��9���9���9E��9+��9���9=��9��9N��9Z��9V��9ɦ�9ӫ�9&��94��95��95��9��9x   x   c��9h��9���9b��9(��9��9"��9���9!��9��9٬�9���9(��9���9���9(��9֫�9v��9*��9_��9���9}��94��9��9��9M��9���9 ��9	��9i��9x   x   ۨ�9���9���9
��9��9]��9ì�99��9w��9���9ث�93��9ة�9k��9���95��9���9��9'��9��9��9ɫ�9_��9��9��9٩�9���9T��9���9ƪ�9x   x   Q��9��9;��9:��9%��9Ƭ�9Ѯ�9U��9���9٨�9k��99��9u��9S��9c��9���9ܨ�9-��9���9;��9@��9���9ī�9J��9��9���9���98��9
��9���9x   x   ��9_��9d��9Ū�9���99��9S��9C��9���9̬�9ѭ�9K��9ܫ�9���9$��9ҫ�9���9��9Ԫ�9���9���9#��9��9���9!��9��9���9Ī�9V��9���9x   x   ��9l��9&��9ë�9"��9v��9���9���9ϫ�9���9���9«�9���9���9׫�9%��9���9	��9ت�9���9@��9n��9��9O��9j��9n��9���9��9���9���9x   x   A��9r��9��9Z��9��9���9٨�9ͬ�9���9��98��9߫�9W��9l��9���9��9���9���9ѩ�9��9���9��9"��9���9a��9��9���9��9ԫ�9o��9x   x   ���9ɬ�9x��9צ�9۬�9׫�9o��9׭�9���90��9	��9��9f��9���9���9��9��9 ��9Ӫ�9��9���9��95��9���9���9���9���9��9��9���9x   x   ��9��9��9G��9���96��95��9I��9���9۫�9��9��9L��9#��9���9ͪ�9���9��9���9���9��9��9W��9��9?��9z��9ë�9��9=��9���9x   x   ��9v��9"��9��9$��9ש�9t��9٫�9���9Z��9h��9I��9-��9A��9���9���9���9ѫ�9«�9֪�9��9���9!��9��9ڧ�9���9H��9+��9��9���9x   x   {��9��9ʦ�9���9���9k��9O��9���9���9k��9��9"��9F��9L��9��9���9ū�9>��9���9��9W��9���9��9s��9���9��9~��9���9]��9��9x   x   4��9_��9`��9���9���9���9c��9(��9ګ�9���9~��9���9���9��9��9Z��9��9���9���9:��9���9���9��9��9o��9#��9���9��9���9h��9x   x   ֨�9���9���9D��9%��99��9���9ԫ�9(��9��9��9˪�9���9���9Y��9x��9��9���9:��9���9��9���9���9b��9*��9W��9m��9X��9��9���9x   x   ���9��9���9,��9׫�9���9ߨ�9ɧ�9���9���9��9��9���9���9��9��9(��9F��9%��9<��9Ѭ�9֬�9ʩ�9���94��9j��9���9t��9ʨ�9E��9x   x   ���9k��9��9���9y��9��9.��9��9	��9���9"��9��9ͫ�98��9���9���9G��9|��9Y��9���9���9��9!��9ƫ�9���9?��9���9Ĩ�95��9���9x   x   ���9���9g��9:��9+��9$��9���9Ϫ�9ت�9̩�9Ӫ�9���9���9���9���9;��9'��9X��9���9~��9���9
��9;��9���9��9ϫ�9��9֪�9>��9���9x   x    ��9[��9���9��9\��9���9>��9���9���9��9��9���9ت�9��9>��9���9>��9���9��9l��9x��9֩�9���9��9���9��9g��9ѫ�9y��9��9x   x   U��9���9���9N��9���9��9<��9���9@��9���9���9��9��9X��9���9��9Ӭ�9���9���9x��9��96��9��9���9���9N��9���9T��9/��9s��9x   x   ���9��9'��9Z��9|��9ƫ�9���9!��9p��9��9��9��9���9���9���9���9׬�9��9��9֩�99��9��9���9(��9���9���9���97��9+��9h��9x   x   ݧ�9���9;��9W��96��9e��9ī�9��9#��9��92��9\��9��9��9��9���9ѩ�9#��9;��9���9��9���9=��9���98��9"��9��9k��9��9���9x   x   ���9���9٨�9Ǧ�9��9��9K��9���9R��9���9���9��9��9x��9��9b��9���9���9���9��9���9'��9���9\��92��9ƫ�9���9ۤ�9���9��9x   x   Ĭ�9��9���9ϫ�9 ��9��9��9!��9n��9b��9���9?��9ܧ�9���9o��9+��95��9���9��9���9���9���95��91��98��9���9��9���9���9>��9x   x   ���9*��9���9'��9O��9ة�9���9��9n��9��9���9y��9���9��9 ��9S��9k��9=��9ͫ�9 ��9I��9���9 ��9ū�9���9\��9��9G��9��9��9x   x   ~��9K��9���90��9���9���9���9��9���9���9���9ǫ�9C��9|��9���9i��9ª�9���9��9e��9���9���9��9���9��9��9���9c��9ά�9.��9x   x   (��9��9���94��9��9T��9=��9���9��9��9��9��9'��9���9��9[��9x��9ƨ�9ת�9ӫ�9Y��92��9k��9ޤ�9���9I��9f��9��9��9	��9x   x   ���9��9`��98��9	��9���9��9R��9«�9ի�9ܥ�9=��9��9^��9���9��9ɨ�98��9<��9w��90��9)��9��9���9���9��9Ϭ�9��9��9���9x   x   ��9���9ϭ�9��9k��9ª�9���9���9���9q��9���9���9���9���9k��9���9C��9���9���9��9r��9g��9���9��9=��9��9/��9��9���9׭�9x   x   Ŧ�9G��9���9]��9���9���9@��9���9w��9c��9p��9ק�9_��9ߧ�9H��9��9��9���9֥�9d��9K��97��9{��9���9x��99��9è�9F��9[��9&��9x   x   B��9u��9��9t��9o��9��94��9��9B��9���9Y��9���9ݦ�9��9���9˥�9��9 ��9F��9��9Q��9���9o��9���9z��9��95��9���9���99��9x   x   ���9��9>��9���9֥�9��9K��9���9H��9���9��9���9��9)��9���9���9���9��9��9���9C��9��9���9ը�9���9��9��9C��9��9��9x   x   _��9r��9���9���9���9M��9���9��9���9���9B��9q��9���9u��9���9p��9 ��9D��9��9��9*��9���9��9��9ۤ�9��9c��9n��9���9!��9x   x   ���9n��9֥�9���9���9æ�9t��9g��9ި�9f��9֣�9���9Ȩ�9���9���9ޥ�9���9%��9���9��9��90��9J��9ث�9���9y��9©�9D��9 ��9ܥ�9x   x   ã�9��9��9N��9¦�96��9���9;��9���9���9m��9m��9��9&��9��9Ψ�9Z��9���9��9K��9d��9��9E��9��9���9���9%��9��9'��9ƥ�9x   x   A��93��9G��9���9s��9���9K��9̧�9���9���9/��94��9��9���9Z��9���9��9]��9Z��9 ��9Ŧ�9Ǩ�9��9æ�98��9H��9Ө�9ܤ�9ԧ�9���9x   x   ���9��9���9��9g��9;��9ϧ�94��9(��9���9���9���9R��9��9S��9��9x��9Y��9$��9J��9¦�9ţ�9Ũ�9֨�9v��9ç�93��9���9��9���9x   x   w��9C��9I��9���9ۨ�9���9���9)��9ש�9��9���9K��9��9���9!��9���9]��9D��9���9���9s��9���9���9r��9���9e��9��9���9���9?��9x   x   d��9���9���9���9e��9���9���9���9��9
��9��9���9���9%��9��9|��9��9Ϩ�9��9���9
��9Q��9���9m��9X��9R��9��9���9̩�9G��9x   x   q��9[��9��9A��9ף�9p��9,��9���9���9��9w��9ר�9��9��9��9��9Ȥ�9a��9k��9��9���97��9���9f��9C��9B��9��9��96��9ƥ�9x   x   ֧�9���9���9o��9���9l��9.��9���9R��9 ��9Ԩ�9���9��9U��9P��9ҥ�9Ԩ�9���9B��9���9Y��9j��9��9��9���9v��9~��9���9��9���9x   x   c��9ܦ�9ާ�9���9Ǩ�9��9��9R��9��9���9��9��9n��9W��9!��9E��9���9Ѧ�9��9���9ç�9Q��9���9h��9c��9ަ�9��9d��9��9l��9x   x   ܧ�9 ��9&��9x��9���9&��9���9��9���9"��9��9X��9W��9Ť�9��9Ȧ�9��9���94��9M��9��9N��9m��9���9z��9̧�9���9u��9���9��9x   x   G��9���9���9���9���9��9X��9R��9��9��9��9P��9!��9��9��9[��9��9��9\��9=��9��9ʤ�9���9ݦ�9��9գ�9Σ�9���9���9���9x   x   ��9˥�9���9p��9ޥ�9Ҩ�9���9��9���9z��9��9ե�9F��9Ʀ�9Z��9ã�9ϧ�9��9���9��9��9+��9��9��9��9���9F��9m��95��9��9x   x   ��9��9���9��9���9X��9��9u��9Z��9��9Ť�9Ҩ�9���9���9��9ϧ�9���9��9���9P��9���9���91��9M��9R��9��9���9b��9���9|��9x   x   ���9!��9��9D��9$��9���9Z��9U��9F��9Ψ�9b��9���9զ�9���9��9��9��9���9ԣ�9��9a��9���9R��9n��9��9 ��9I��9��9��9���9x   x   ץ�9E��9��9��9���9��9Y��9$��9���9��9m��9?��9��95��9Z��9���9���9ӣ�9���9���9���9R��9���9���9���9^��9���9!��9��9��9x   x   b��9��9���9��9��9L��9��9L��9���9���9��9���9���9J��99��9��9L��9��9���9Ū�9��9���9��9l��9)��9��9p��9D��9���9���9x   x   J��9L��9C��9+��9��9`��9Ǧ�9���9s��9��9���9X��9���9��9��9��9���9a��9���9��9p��9���9��9���9���9���9��9���9g��9z��9x   x   5��9���9��9���93��9��9ʨ�9ţ�9���9O��9<��9j��9R��9Q��9ʤ�9/��9���9���9W��9���9���9m��9���9r��9R��9'��9[��9��99��9���9x   x   z��9k��9���9��9J��9A��9��9¨�9���9���9���9��9���9m��9��9��9+��9S��9���9��9��9���9'��9r��9j��9��9���9=��9S��9Ŧ�9x   x   ��9���9֨�9��9ث�9��9æ�9Ҩ�9s��9i��9j��9��9i��9���9٦�9!��9M��9o��9���9l��9���9u��9r��9��9���9w��93��9ʩ�9%��9X��9x   x   y��9y��9���9ޤ�9��9���98��9s��9���9U��9D��9���9d��9v��9��9��9O��9��9���9)��9���9Q��9j��9���9���9l��9ޤ�9���9_��9��9x   x   ;��9��9��9��9v��9���9J��9ħ�9g��9O��9E��9u��9��9Χ�9أ�9���9��9��9`��9��9���9+��9��9x��9s��9`��9���9L��9��9$��9x   x   Ȩ�95��9��9e��9ũ�9'��9֨�95��9��9��9��9~��9��9���9̣�9G��9���9E��9���9o��9��9Y��9���90��9ߤ�9���9s��9F��9��9��9x   x   I��9���9D��9q��9H��9��9ܤ�9���9���9���9��9���9d��9t��9��9k��9b��9��9��9D��9���9ߦ�9B��9Ʃ�9��9H��9B��9���9��9���9x   x   Y��9���9��9���9���9#��9ا�9��9���9˩�99��9��9��9���9���95��9��9��9��9æ�9j��9:��9S��9)��9`��9��9��9��9���9է�9x   x   !��9;��9���9 ��9��9ƥ�9���9���9>��9F��9ƥ�9���9f��9��9���9��9{��9���9��9���9}��9���9Ħ�9V��9��9%��9��9���9٧�9���9x   x   [��9��9ê�9'��9٣�9ا�9���9c��9���9:��9���9W��9���9ߤ�9S��9	��9��9���9^��9���9��9ӥ�9s��9֤�9��9��9���9���9ި�9���9x   x   ��9H��9���9���9Ƣ�9,��9���9u��9���9��9\��9ѧ�9���9ģ�9E��9���9>��9���9��9)��9^��9���9+��9آ�9���9F��9���9��9ܦ�9���9x   x   ª�9���9Z��9��9���9ѥ�9i��9���9��9"��9@��9U��9ܢ�9k��9D��9��9|��99��9���9s��9Ѧ�9���9��9���9ۦ�9w��9���9 ��9���97��9x   x   ,��9���9��9���99��9���9"��9Ԩ�9���9��9��9��9��9��9���9R��9f��9>��9��9���9>��9��9b��9`��9Ԧ�9/��9��9J��9��9L��9x   x   ڣ�9Ƣ�9���96��9w��9=��9��9p��9���9���9ˤ�9��9���9e��9���9��9B��9���9��9���9���9i��9y��9ʤ�9ߦ�9á�9���9���9���9���9x   x   ֧�9+��9ѥ�9���9;��9��9{��9��9g��9���9)��9���95��9R��9���9m��9��9��9��9$��9'��9L��9#��9C��9���9���9���93��9Х�9ɦ�9x   x   ���9���9k��9$��9��9x��9N��9��9.��9��9!��9*��9���9��9��9Ӥ�9��9��9���9ħ�9P��9���9���9���9���9���9O��9¥�9���9���9x   x   _��9v��9���9Ө�9p��9���9��99��9
��9���9��9>��9I��9[��9���9Ҥ�9��9���9���9���9��9��9���9֤�9]��9���9^��9���9>��92��9x   x   ���9���9��9���9���9f��9+��9��9v��9ا�9˦�9��9���9§�9֢�9��9���9Ȥ�9£�9v��9��9���9��9���9���9���9ҥ�9���9ޤ�9��9x   x   8��9��9 ��9��9���9���9��9���9ק�9���9'��9d��9���9���9���9Ȥ�9���9���9��9���9���9���9��9��9{��9P��94��9^��9���9]��9x   x   ���9\��9@��9��9Ȥ�9+��9!��9��9Ȧ�9$��9F��9��9��9��9a��9n��9˥�9���9ۧ�9ͩ�9N��9٤�9���9"��9l��9W��9���9ר�9���9 ��9x   x   X��9ϧ�9U��9��9��9���9,��9<��9��9`��9��9��90��9��9M��9���9N��9���9��9���9j��9���9ţ�9)��9!��9���9`��9��9��9O��9x   x   ���9���9��9��9���96��9���9F��9���9���9��9/��9��9F��9?��9��9U��9X��9ϧ�9���9y��9!��9���9)��9���9>��9֥�9r��9)��97��9x   x   ۤ�9ȣ�9j��9��9b��9K��9��9\��9Ƨ�9���9��9��9A��9���9ܤ�9���9��9���9���9w��9$��9l��9:��9��9���9��9^��9��9��9Υ�9x   x   Q��9I��9F��9���9���9���9��9���9ܢ�9��9a��9K��9?��9ߤ�9���9���9���9z��9t��9.��9��9��9���91��9`��9���9���9M��9���9��9x   x   
��9���9��9Q��9ޤ�9o��9Ӥ�9Ԥ�9��9Ǥ�9m��9���9��9���9���9$��9(��9��9J��9���9���9p��9ݩ�9���9+��9f��9��9d��9���9���9x   x   ��9<��9~��9h��9@��9��9��9~��9��9���9˥�9N��9Q��9 ��9��9&��9��9��9e��9q��9���9���9L��9���9���9פ�9���9��9z��9}��9x   x   ���9���99��9A��9���9��9
��9���9Ȥ�9���9���9���9W��9���9y��9��9��9"��9��98��9���9���9��9۪�9e��9Ʃ�9˥�9-��9p��9#��9x   x   \��9��9���9��9��9��9���9���9���9��9٧�9��9ϧ�9���9t��9K��9e��9���9���9*��9��9+��9��9���9I��9O��9,��9���9���9T��9x   x   ���9*��9u��9���9���9��9§�9���9t��9���9Щ�9���9���9{��9/��9���9p��9<��9'��9���9.��9d��9���9��9���9a��9A��9V��9G��9ҥ�9x   x   ��9`��9Ϧ�9;��9���9)��9T��9��9��9���9Q��9f��9~��9%��9��9���9|��9���9��9(��9���9��9���9��9؟�9U��9;��9��9	��9���9x   x   ҥ�9���9���9��9k��9N��9���9��9���9���9դ�9���9"��9j��9��9m��9���9���9)��9`��9��9k��9��9p��9b��9���9��9q��9-��9ѥ�9x   x   s��9+��9��9`��9w��9��9��9���9	��9��9���9���9���99��9���9ߩ�9H��9��9��9���9���9��9���9թ�9P��9��9 ��9���9��9��9x   x   դ�9ڢ�9���9`��9ͤ�9E��9���9ؤ�9���9��9%��9'��9-��9��99��9���9���9��9���9��9���9n��9֩�9B��9o��9w��9��9R��9)��93��9x   x   ��9���9ۦ�9Ҧ�9ߦ�9���9���9^��9���9|��9m��9!��9���9���9a��9&��9���9h��9E��9���9ٟ�9_��9R��9r��9���9��9���90��9���9}��9x   x   }��9G��9y��9.��9ġ�9���9���9���9���9O��9Y��9���9=��9��9���9c��9Ф�9ȩ�9K��9[��9T��9���9��9s��9��9^��92��9���92��9i��9x   x   ���9���9���9���9���9���9N��9\��9ϥ�92��9���9\��9֥�9^��9���9��9���9ҥ�9+��9C��9=��9��9!��9��9���92��9=��9���9ȥ�9���9x   x   ���9��9��9G��9���95��9¥�9���9���9b��9ب�9��9t��9��9L��9f��9��9-��9���9V��9��9p��9���9T��91��9���9���9��98��9=��9x   x   ��9ަ�9���9��9���9ѥ�9���9A��9ݤ�9���9���9��9,��9��9���9���9y��9r��9���9F��9	��9+��9��9(��9���95��9ʥ�96��9ԣ�9t��9x   x   ���9���9>��9N��9���9ʦ�9���92��9��9\��9��9M��98��9ͥ�9��9���9y��9#��9V��9ѥ�9���9֥�9��9-��9{��9f��9���9=��9s��9��9x   x   ��9���9=��9���9���99��9��9r��9��9w��9��9y��9��9���9���9+��9���9���90��9���9���9W��9��90��9n��9���9���9���9��9��9x   x   ��9��9a��9P��9ˣ�9���9���9���9g��9>��9��9���9��9ܧ�91��9@��9+��9��9^��9��9��9ã�9���9���9}��9a��9���9���9��9z��9x   x   <��9a��9���9ǧ�9���9(��9ۧ�9z��94��96��9/��9q��9A��9��9	��9��9ۥ�9ǥ�9<��9y��9��9&��9E��9��9���9/��9Ԧ�9N��9���9$��9x   x   ��9N��9Ƨ�9���9;��9���9��9��9|��9���9���9���9���9���9[��9]��9ؤ�9���95��9x��9V��9פ�9���9���9?��9٧�9ؤ�9ĥ�9ǥ�9f��9x   x   ���9Σ�9���99��9���9���9G��9��9���9��9��9��9���9���9���9��9���9��9c��9���9���9���9ҩ�9���9.��9��9���9���9��9���9x   x   6��9���9'��9���9���9���9;��9��9��9���9~��9��9,��9k��9j��9(��9��9 ��9��9��9e��9���9��9��9��9��9æ�9b��9��9
��9x   x   ��9���9ڧ�9
��9L��9?��9��9��9��9���9g��9��9&��9G��9Y��9P��9=��9���9���9f��9g��9]��9$��9֥�9G��9���9���9P��9��9���9x   x   r��9���9z��9��9��9��9��9~��9ӥ�9��9å�9N��9���9٤�9��9��9���92��9^��9���9ӡ�9O��9@��9;��9:��9���9I��9���9���9���9x   x   ��9i��96��9x��9���9��9��9ե�9ȥ�9���9���9��9%��9���9��9���9��9A��9���9`��9f��9���9e��9���9���9`��9���9���9���9��9x   x   t��9?��98��9���9��9���9���9��9���9k��9Ӧ�9��9���9���9 ��9ץ�9z��9
��9+��9d��9��9��9���9U��9���9���9Y��9N��9��9���9x   x   ��9��9/��9���9��9��9f��9¥�9���9Ԧ�9'��9צ�9<��9���9"��9��9l��9g��9Ѥ�9���9y��9k��9Σ�9���9���9'��9���9t��9���9Q��9x   x   x��9 ��9m��9 ��9��9��9��9P��9��9��9ަ�9��9ߤ�9���9x��9X��9��9���9P��9���9���9k��9���9���9*��9է�9j��9ĥ�9c��9��9x   x   ��9��9:��9���9���9(��9"��9���9(��9���9>��9ߤ�9��9��9Z��9��9��9§�9���9���9r��9 ��9٦�9��9ؤ�9p��9��9ާ�9x��9���9x   x   ���9ާ�9��9���9���9m��9H��9ؤ�9���9���9���9���9��9;��9D��9���9��9���9O��9���9���9^��9|��9S��9b��9:��9H��9���9���9��9x   x   ���9+��9��9\��9���9m��9Y��9��9��9 ��9#��9{��9Z��9E��9m��9���9ǣ�9��9&��9���9���9%��9N��9Υ�9��9��9��9'��9���9#��9x   x   .��9<��9~��9Z��9��9'��9T��9��9���9إ�9��9V��9���9���9���9���9���9n��9���9���9,��9g��9���9���9��9~��9��9���9j��9(��9x   x   ��9*��9٥�9٤�9���9��9<��9���9��9y��9l��9��9��9��9ʣ�9���9���9$��9 ��9ɤ�9
��9���9B��9A��9���9m��9���94��9.��9+��9x   x   ���9���9ƥ�9���9��9���9���9/��9:��9��9e��9���9ŧ�9���9��9n��9$��9��9���9��9ŧ�9���9��9��9���9���9ˤ�9���9ܧ�9���9x   x   0��9c��9<��94��9d��9��9���9^��9���9-��9Ѥ�9P��9���9O��9'��9���9���9���9n��9U��9$��9���9���9 ��9C��9���9Ȧ�9��9���9V��9x   x   ��9��9y��9y��9���9��9d��9���9d��9a��9���9���9��9���9���9���9̤�9z��9X��9���9��9���9J��9 ��9ԥ�9ޣ�98��9���9���9@��9x   x   ���9 ��9��9W��9���9e��9c��9ס�9e��9	��9y��9���9n��9���9���9/��9��9���9)��9��9���9%��9���9���9���9e��9��91��9]��9���9x   x   Z��9���9%��9פ�9���9���9Z��9K��9���9	��9j��9p��9��9]��9)��9f��9���9���9���9���9)��9p��9���9#��9���9f��9£�9Ѩ�9��9��9x   x   ��9���9C��9���9֩�9���9#��9<��9e��9���9̣�9���9ئ�9|��9P��9���9D��9��9���9K��9���9���9��9I��9���9��9ץ�9���9ޤ�9H��9x   x   3��9���9��9���9���9��9֥�9?��9���9R��9���9���9��9R��9ʥ�9��9B��9��9���9��9���9#��9I��9���9)��93��9"��9��9��9���9x   x   j��9}��9���9;��9-��9��9D��99��9���9���9���9+��9֤�9b��9��9��9���9���9G��9ۥ�9���9���9���9)��9���9w��9���9ɧ�9���9���9x   x   ���9e��9.��9ا�9 ��9��9���9���9b��9���9%��9է�9p��98��9��9���9o��9���9���9ޣ�9d��9d��9��95��9w��9^��9W��98��9i��9,��9x   x   ���9���9֦�9ؤ�9���9æ�9���9J��9���9X��9���9r��9��9G��9��9��9���9ͤ�9Ȧ�97��9��9ã�9إ�9'��9���9R��9���9��9���9&��9x   x   ���9���9P��9ȥ�9���9b��9Q��9���9���9M��9s��9ǥ�9ߧ�9���9'��9���9/��9���9��9���93��9Ѩ�9���9��9ȧ�96��9��9{��9���9���9x   x   ��9ޢ�9���9ĥ�9��9��9��9���9���9 ��9���9e��9t��9���9���9n��90��9ݧ�9���9���9^��9��9ۤ�9��9���9e��9���9���9]��9��9x   x   ��9z��9$��9d��9���9��9���9���9��9���9R��9��9���9��9#��9+��9/��9���9U��9D��9���9��9J��9���9���9,��9'��9���9��9��9x   x   ���9���9���9Ţ�9r��9*��9���9���9_��9���9Ϧ�9p��9+��9���9ǩ�9ߤ�9���9i��9��9���9e��91��9���9Ч�9զ�9���9
��9w��9֤�9���9x   x   ��9���9l��9|��9���9ң�9���9���9Y��9���9��9F��9$��9��9B��9ڥ�9D��9���9���9��9��9M��9@��9)��9N��9��9��9��9���9���9x   x   ���9s��9U��9*��9���9]��9��9��9���9���9���9���9��9w��9զ�9O��9���9���9��9���9��9Ң�9٢�9��9٧�9C��9���9Ĩ�9���90��9x   x   â�9��9%��9��9���9��9��9ħ�9���9���9��9���9���97��9��9���9t��9W��9���9���9Y��9���9���9[��9���9á�9���9���9s��9��9x   x   v��9���9���9���9$��9W��9���9���9Ф�9���9���9.��9&��9g��9e��95��9���9���9ݤ�9��9���9��9���9̩�9���9'��9��9f��9���9���9x   x   /��9У�9`��9��9U��9���9p��9Q��9��9N��9ɤ�9���9^��9D��9,��9���9���9ʥ�9ʢ�9g��9Χ�9���9��9���9��9��9}��9���9	��9���9x   x   ���9���9 ��9��9���9n��9@��96��9���9T��9Ƥ�9x��9���9��9Q��9ͦ�9Ȩ�9���9W��9k��9A��9ӧ�9���9��9��9��9;��9u��9<��9ڦ�9x   x   ���9���9��9ŧ�9���9O��97��90��9\��9ǣ�9x��9���9���9���94��9r��9���9{��9��9���9ק�9^��9J��9���9i��9{��9��9��9ͩ�91��9x   x   _��9V��9���9���9Ԥ�9��9���9\��9̤�9���95��9���9o��9W��9���9��9y��9ޥ�9���9���9��9t��9���9���92��9"��9��9Ĥ�9I��9��9x   x   ���9���9���9���9���9P��9T��9ƣ�9���9���9���9���9r��9w��9\��9���9��9#��9���91��9���9Ц�9��9��9���9��9@��9���9���9a��9x   x   Ѧ�9��9���9��9���9Ȥ�9Ȥ�9v��94��9���9X��9���9���9��9��9c��9B��9Q��9���9I��9���9���9���9b��9Ф�9}��9��9n��9v��9���9x   x   q��9G��9���9���9.��9���9{��9���9���9���9���9B��9y��9U��9���9ϧ�9��9��9z��9b��9ܤ�9a��9K��9���9���9c��9���9��9���9f��9x   x   ,��9#��9��9���9%��9a��9���9���9n��9n��9���9{��9��9Z��9?��9��9ۤ�9���9���9���9¤�9i��9��9'��90��9��9V��9E��9��9��9x   x   ���9��9~��94��9e��9H��9��9���9[��9z��9��9R��9[��9f��9��9���9���9��9��9v��9 ��9���9��9w��9��9~��9���9��9ߤ�9l��9x   x   ȩ�9B��9צ�9��9a��9*��9P��96��9���9a��9��9���9=��9��9v��9���9���9���9	��9��9��9���9��9��9L��9��9���9���9C��9���9x   x   ��9إ�9S��9 ��97��9���9ͦ�9q��9��9���9c��9ҧ�9��9���9���9��9���9��9��9���9���9��9\��9f��9|��9���9���9���9���9���9x   x   ���9E��9���9u��9���9��9ƨ�9���9z��9 ��9B��9��9ݤ�9���9���9���9֤�9~��9��9���9���9ĥ�9���9L��9<��9��9^��9u��9
��9Ť�9x   x   h��9���9���9T��9���9ϥ�9���9}��9��9%��9M��9ߩ�9���9��9���9��9���9���9��9o��9���9��9P��97��9���9(��9Y��9��9q��9��9x   x   ��9���9$��9���9ޤ�9ɢ�9U��9��9���9���9���9y��9���9��9��9��9���9��9��9���9&��9���9���93��9-��9���9<��9���9ɣ�91��9x   x   ���9��9���9���9���9f��9j��9��9���93��9L��9_��9ª�9x��9��9���9���9p��9���9��9e��9`��9���9E��9���9���9X��9��9��9é�9x   x   d��9��9��9Y��9���9ԧ�9@��9ا�9��9���9���9��9���9��9��9���9���9���9(��9c��9���9���9g��9/��9W��9/��9a��9	��9D��9	��9x   x   2��9K��9Ԣ�9���9��9���9է�9`��9v��9ͦ�9��9a��9h��9���9���9��9å�9��9���9X��9���9��9���9���9���9��9���9*��9���9���9x   x   ���9?��9֢�9���9���9��9���9I��9���9��9���9I��9��9��9��9`��9���9S��9���9���9l��9���9���9��9*��9��9ݢ�99��9f��9���9x   x   ԧ�9+��9��9Y��9ũ�9���9��9���9���9��9c��9���9%��9x��9��9h��9K��95��99��9D��91��9å�9
��9���9��9ƥ�9m��9"��9���9��9x   x   Ԧ�9N��9ۧ�9���9���9	��9��9i��94��9���9Ϥ�9���91��9��9L��9y��9<��9���91��9���9O��9���9)��9��9W��9���9أ�9?��9ע�9���9x   x   ���9��9A��9ơ�9#��9��9
��9|��9��9��9}��9d��9��9���9��9���9���9!��9���9Ħ�9/��9��9��9ƥ�9���9��9&��9���9@��9b��9x   x   ��9��9���9���9��9~��9=��9��9��9D��9��9���9S��9���9���9���9d��9X��9<��9Y��9a��9���9ڢ�9l��9أ�9+��9���9t��9��9Z��9x   x   z��9��9Ĩ�9ţ�9g��9���9t��9���9ä�9���9k��9��9D��9��9���9���9y��9	��9���9��9	��9*��98��9��9A��9���9q��9���9���9��9x   x   դ�9���9���9q��9���9
��9=��9Ω�9H��9���9w��9���9��9ߤ�9D��9���9��9l��9̣�9��9C��9��9h��9��9֢�9@��9��9���9��9��9x   x   ��9���91��9��9���9���9ݦ�91��9���9a��9���9f��9��9m��9��9��9Ƥ�9��90��9���9��9���9���9��9���9c��9[��9��9��9[��9x   x   n��9U��9G��9#��9դ�9���9<��9���9g��9U��9���9z��9t��9J��9$��9��9��9a��9>��9��9��9S��9^��9y��9���9Z��9���9˪�9���9f��9x   x   W��9���9ŧ�9���9	��9��9���9?��9e��9Y��9���9i��9|��9F��9'��9��9��9>��9S��9��9Ƨ�9���9g��9��9���9���9��9��9���9��9x   x   F��9ħ�9��9���9i��9���9���9��9R��9{��9ǧ�9���9X��9���9���9ب�9��9c��9���9ɩ�93��9?��9���9O��9.��9p��9���9N��9=��9ͦ�9x   x   "��9~��9���9/��9���9���9���9���9��9���9��96��9���9���9ͦ�9e��9���9/��9K��9L��9��9��9P��9ۧ�9+��9ê�9ӥ�9��9��9���9x   x   Ԥ�9	��9k��9���9���9��9=��9/��9.��9���9��9���9���9	��9=��9��91��9���9���9[��9���9d��9��9���9���9)��9��9��9h��9p��9x   x   ���9��9���9���9��9��9a��9���9��9-��9֨�9���9=��9���9���9���9��9���9��9G��9 ��9Ҫ�9l��9���9���9Ω�9���9��9	��9y��9x   x   =��9���9���9���9<��9b��9��9��9Ϧ�9o��9c��9���9���9���9ʩ�9Ч�9���9|��9s��90��9���9A��9թ�9���98��9f��9���94��9��9��9x   x   ��9?��9��9���91��9���9��9���9��9{��9���9��9���9���9Z��9���9���9$��9n��9ީ�9���9ª�9>��9��9��9���9���9^��9z��9���9x   x   e��9e��9Q��9��9.��9��9Φ�9��9���9ŧ�9v��9|��9S��9���9Q��9k��9=��9ƨ�9���9"��9��9H��9
��9Ы�9��9̨�9���91��9���9e��9x   x   V��9Z��9|��9���9���9.��9o��9{��9Ƨ�9y��9��9���9���9n��9r��9���9���9���9B��9v��9��9���9W��9���9<��9��9��9l��9ʦ�9���9x   x   ���9���9ʧ�9��9}��9ը�9e��9���9v��9��9��9���9{��9\��9x��9R��9���9)��9��9���9:��9.��9;��9��9���9���9٨�9٩�9���9���9x   x   z��9e��9���95��9���9���9���9��9|��9���9���9���9���9���97��9��9_��9ͦ�9*��9��9Ѧ�9���9ƨ�9���9���9ڧ�9k��96��9l��9��9x   x   t��9|��9Y��9���9���9:��9���9���9S��9 ��9z��9���9m��9G��9���9,��9`��9P��9=��96��9-��9��9Ҫ�9u��9���9���9���9u��9V��93��9x   x   K��9E��9���9���9
��9���9���9���9���9m��9Z��9���9G��9���9)��9.��9���9���9��9���9*��9ԩ�9|��9>��9���9p��9���9���9;��9���9x   x   $��9$��9���9Ϧ�9@��9���9̩�9X��9O��9o��9z��97��9���9,��9Ũ�9;��9	��9ݧ�9[��9w��9��9w��9���9?��9U��9>��9���9>��9��9��9x   x   ���9��9Ԩ�9c��9��9���9Χ�9���9l��9���9V��9��9*��9.��99��9ѩ�9���9ۥ�9-��9���9=��9��9���9n��9x��9T��9n��9 ��9���9���9x   x   ��9��9��9���9/��9��9���9���9@��9���9���9`��9]��9���9
��9���9=��9��9���9Ч�9���9��9��9-��93��9ѧ�9a��9��9��9e��9x   x   _��9@��9h��92��9���9���9|��9!��9Ĩ�9���9-��9Φ�9O��9���9��9ܥ�9��9���9���9a��9K��9N��9��9���9��9���9ا�9
��9��9���9x   x   @��9P��9���9N��9���9��9u��9n��9���9E��9��9,��9@��9��9Z��90��9���9���9���9D��9:��9���9y��9���9h��9���95��9���9��9m��9x   x   ��9 ��9ǩ�9N��9`��9F��9/��9��9%��9t��9���9��96��9���9v��9���9̧�9`��9?��9��9���9p��9���9w��9���9���9��9-��9'��9��9x   x   ��9ȧ�92��9��9���9 ��9���9���9��9��9>��9Ϧ�9,��9(��9��9?��9���9M��95��9���9���9Ҩ�9*��9���9���9*��9���9"��9���9Ĩ�9x   x   P��9���9?��9��9b��9Ϫ�9@��9���9H��9��9-��9���9��9ѩ�9x��9��9��9V��9���9t��9ը�9H��9���9Ѩ�9��9���9���9"��9y��9e��9x   x   ^��9g��9��9P��9��9k��9ԩ�9@��9��9Y��9:��9Ũ�9Ԫ�9|��9���9���9ۣ�9��9t��9���9)��9���9���9/��9��9��9��9���9���9ק�9x   x   s��9��9P��9٧�9���9���9��9��9̫�9���9��9���9w��9=��9@��9q��9+��9���9���9y��9���9Ҩ�9/��9���9���9���9i��9Y��9Y��9��9x   x   ���9���9.��9(��9���9���99��9��9ߧ�9;��9���9���9���9���9S��9x��94��9��9g��9���9���9��9��9���96��9��9���9.��99��9���9x   x   X��9���9r��9���9*��9Ω�9c��9���9Ϩ�9��9���9ۧ�9���9p��9=��9U��9Ч�9���9���9���9*��9���9��9���9��9Ы�9&��9��9:��9_��9x   x   ���9���9���9إ�9��9���9���9���9��9��9ۨ�9l��9���9���9���9n��9`��9է�90��9
��9���9���9��9j��9���9$��9���9���9��9���9x   x   ɪ�9��9K��9
��9z��9��93��9_��90��9l��9ک�96��9w��9��9=��9��9��9��9���9*��9"��9#��9���9Z��9-��9}��9���9��9���97��9x   x   ���9���9?��9��9l��9
��9��9z��9���9ɦ�9���9f��9[��99��9��9���9��9��9��9'��9���9v��9���9\��97��9?��9��9���9��9���9x   x   b��9��9˦�9���9l��9z��9��9���9c��9���9���9��95��9���9��9���9h��9~��9l��9���9Ȩ�9d��9ק�9��9���9]��9���98��9���9j��9x   x   ���9ޫ�9u��9��9��97��9d��9���9A��9l��9k��9ũ�9w��9��9b��9y��9��9��91��9`��9��9U��9@��9L��9��9��9��9ŭ�9���9��9x   x   ݫ�9���9b��9��9��9���9���9���9���9���9���9ߪ�9���9&��9���9ӫ�9ê�9Q��9��9T��9��9��9���9��9B��9��9��9���9���9���9x   x   t��9b��9���9p��9���9F��9���93��9��9z��9���9���9���9'��9y��9W��9���9o��9Ѫ�9ͬ�9���9���9ά�9̫�9���9c��9ݬ�9��9M��9���9x   x   ��9��9r��9%��9��9���9=��9.��9{��99��9��9��9ԫ�9���9M��9G��9���9:��9���9ث�9|��9���9?��9���9��9���9J��9	��91��9���9x   x   ��9��9���9{��9��9	��9f��9���9t��9��9b��9S��9Z��9��9��9y��9+��9$��9��9��9̨�9j��9���9���9ڪ�9'��9U��9b��9X��9X��9x   x   5��9���9G��9���9��9���9m��9(��9���9���9`��92��9X��9���9ө�9��9���9��9c��9A��9���9���94��9���9f��9s��9��9��9$��9���9x   x   f��9���9���9;��9g��9n��9���9��9Ȫ�9i��9"��9e��9���9��9���9Ī�9���9���9+��9��9���9��9���9��9i��9���9ܨ�9���9��9j��9x   x   ���9���95��9.��9���9)��9��9ӭ�9��9���9���9���9���9i��9~��9��9���9��9!��9{��91��9���9���9��9ժ�9��9���9L��9���9���9x   x   A��9���9��9z��9s��9���9Ȫ�9��9>��9��94��9���9��9>��9
��9���9k��9"��9̪�9���9���9���9۬�94��9���9 ��9ɫ�9o��9O��9ݮ�9x   x   m��9���9{��98��9��9���9g��9���9��9��9���9~��9i��99��9���9R��9&��9v��9��9���9N��9���9��9(��9��9Ʃ�9��9a��9q��9���9x   x   h��9���9���9��9b��9a��9#��9���94��9���9ͭ�9ȫ�9#��9>��9z��9Ҭ�9֫�9G��9��9��9��9ܯ�9���9���9���99��9ݫ�9���9d��9P��9x   x   ȩ�9ܪ�9���9��9U��9/��9e��9���9���9��9ȫ�9ު�9��9֪�9_��9���94��9ܪ�9���9`��9���9��9���9(��9���9��9���9���9���9���9x   x   y��9���9���9ҫ�9]��9W��9���9���9��9j��9#��9��9���9Z��9x��9��9̫�9j��96��9.��9��9���9ƭ�9ث�9T��9��9���9խ�9��9D��9x   x   	��9%��9(��9���9��9���9��9i��9<��9:��9>��9֪�9\��9���9���9���9O��9���9~��9���9"��9j��9���9j��9��9���9O��9 ��9Y��9ܫ�9x   x   d��9���9{��9P��9��9ѩ�9���9~��9	��9���9|��9_��9w��9���9���9ޫ�9h��9ڪ�9���9��9���9ǫ�9���9��9R��9���9W��9���9���9���9x   x   |��9ԫ�9U��9F��9z��9��9���9��9���9P��9Ѭ�9���9��9���9ݫ�95��9��9��9+��9���9��9Ҭ�9���9w��9`��95��9���9��9���9���9x   x   ��9Ū�9���9���9*��9���9���9���9k��9'��9ҫ�96��9˫�9R��9i��9��95��9l��9X��9��9���9���9Y��9��9G��9��9֫�9r��9��9���9x   x   ��9R��9r��9;��9#��9��9���9��9!��9v��9H��9ު�9i��9���9ܪ�9��9h��9���9���9���9���9ī�9a��9L��93��9Y��9&��9���9��9���9x   x   4��9ު�9̪�9��9��9b��9/��9"��9˪�9��9��9���99��9}��9���9-��9V��9���9>��9���9���9~��9Ů�9&��9���9^��9���9���9��9��9x   x   c��9U��9̬�9٫�9��9@��9��9}��9���9��9߭�9]��9,��9���9��9���9��9���9���9Ω�97��9��9���9���9���9߫�9B��9���94��9���9x   x   ��9��9��9{��9Ϩ�9���9���90��9���9P��9��9���9��9"��9���9��9���9���9���9=��9���9n��9s��9[��9���9���9,��97��9p��9���9x   x   R��9��9���9���9k��9���9��9���9���9���9ܯ�9��9���9g��9ɫ�9լ�9���9ɫ�9|��9��9o��9��9��9���9��9��96��9���9���9"��9x   x   C��9���9ͬ�9?��9���94��9���9���9ݬ�9��9���9���9ǭ�9���9���9���9S��9a��9®�9���9q��9��9{��9A��9Ϋ�9e��9&��9Ϊ�9���9|��9x   x   I��9��9ʫ�9���9���9���9
��9��93��9%��9���9'��9٫�9h��9��9{��9��9P��9%��9���9b��9���9A��9��9���9A��9���9��9���9Q��9x   x   ��9B��9���9���9ت�9f��9i��9ڪ�9���9��9���9���9T��9��9P��9a��9I��92��9���9��9���9��9ѫ�9���9��9��9���9��9��9��9x   x   ��9��9c��9���9'��9r��9���9��9��9ũ�9;��9��9��9���9���96��9��9]��9c��9��9���9��9d��9A��9��9<��9Ҫ�9���9{��9���9x   x   ��9��9ެ�9O��9T��9��9ި�9���9ɫ�9|��9ݫ�9���9���9K��9Z��9���9ԫ�9"��9���9A��90��95��9&��9���9���9Ъ�9٪�9���9��9:��9x   x   ­�9���9��9��9_��9��9���9L��9q��9`��9���9���9٭�9���9���9���9p��9���9���9���97��9���9Ϊ�9��9��9���9���9��9���9��9x   x   ���9���9M��93��9X��9$��9��9���9Q��9o��9f��9���9��9U��9���9���9��9
��9��92��9n��9���9���9���9��9���9��9���9���9̫�9x   x   ��9���9���9���9T��9���9g��9���9ܮ�9���9T��9���9F��9ݫ�9���9��9���9���9��9���9���9"��9z��9P��9|��9���9<��9��9ʫ�9I��9x   x   ��9��9o��9t��9��9ǯ�9ޱ�9ױ�9ð�9���9S��9��9V��9,��9���9|��9���9���9��9/��9���9���9*��90��9/��9+��9���9+��9C��9ݱ�9x   x   ��9t��9 ��9*��9��9���9*��9��9���9���9���9i��9��9w��9&��9��9���9���9��9q��9��9���9m��9ڱ�9��9��9���9̲�9p��9���9x   x   o��9��9֬�9Ȭ�9��95��9��9���9^��9q��9O��9���9���9u��9��9��9���9N��9ͱ�9N��9ɯ�9���9���9Ư�9G��9���9��9M��9���92��9x   x   q��9+��9���9���9��9��9���9x��9w��99��9$��9)��9*��90��9Ա�9���9���9���9#��9���9���9���9��9ڳ�95��9y��9���9v��9���9%��9x   x   !��9��9��9��9s��9��9��9=��9ͯ�97��9��9���9��9���9h��9���9E��9O��9ͯ�9ް�9��9k��9,��9o��9��9I��9���9
��9ͳ�9E��9x   x   ˯�9���99��9��9��9���9���9k��9���9���9˯�9l��9���9���9ڲ�9���9±�9��9���9װ�9Y��9=��9��9~��9���9ˮ�9A��9���9N��90��9x   x   ޱ�9%��9��9���9���9���9��9ұ�9ڲ�9W��9*��9g��9\��9���9ԯ�9ΰ�9��9���9��9���9b��9��9���9x��9x��9���9���9O��9l��9���9x   x   ܱ�9��9���9z��9<��9h��9б�9���9-��9���9���9{��9��9��9@��9U��9ΰ�9߱�9l��9���9���9��9���9��9Q��9���9?��91��9��9��9x   x   ���9���9^��9{��9ѯ�9���9ز�9.��9ˮ�9l��9���9a��9Գ�9A��9���9��9��9Ű�9���9���9˯�9��9հ�9L��9��9
��9)��9ů�9ݭ�9v��9x   x   ���9���9p��9:��96��9���9W��9��9o��9n��9F��9]��9A��9}��9G��9L��9k��9��9��9®�9���9���9���9��9���9а�9β�9Ѱ�9��9���9x   x   T��9���9N��9%��9��9̯�9,��9���9���9D��9��9L��9��9���9��9K��9���9���93��9��9$��9���9k��9İ�9+��9��9`��9���9B��9K��9x   x   ��9k��9���9,��9���9k��9i��9y��9`��9X��9L��9'��9P��9��99��9t��9u��9���9���9��9˯�9���9W��9[��9	��9���9W��9��9b��9��9x   x   V��9��9���9)��9��9���9[��9��9Գ�9>��9��9Q��9��9���9��9���9���9��9ٯ�9´�9`��9���9��9���9b��9<��9���9*��9���9,��9x   x   (��9x��9z��9,��9���9���9���9��9C��9~��9���9��9���9���9ޱ�9���9گ�9n��9���9i��9f��9���9ر�9
��9���9;��9���9���9���9���9x   x   ���9$��9��9ϱ�9c��9ٲ�9ԯ�9D��9���9L��9��96��9��9ݱ�9հ�9���9س�9���9���9��9ϳ�9���9��9԰�95��9|��9_��9���95��9U��9x   x   ��9 ��9��9���9���9���9ϰ�9U��9��9J��9K��9x��9���9���9���9`��9a��9��9ʯ�9���9s��9&��9���9լ�9���9���9���9[��9m��9֮�9x   x   ���9���9���9���9F��9���9��9Ѱ�9��9l��9���9v��9���9گ�9س�9^��9���9[��9���9t��9��9���9]��9d��9p��9���9E��9m��9׮�9_��9x   x   ���9���9K��9���9P��9��9���9��9Ȱ�9��9���9���9��9n��9���9��9_��9���9��9���99��9g��9���9���9��9(��9��9��9j��9���9x   x   ޯ�9��9ұ�9"��9ί�9���9��9o��9���9��9:��9���9د�9���9���9̯�9���9��9���9Ʋ�9���9H��9��9O��9ǲ�9��9	��9"��9J��9ٮ�9x   x   /��9p��9O��9���9ڰ�9ְ�9���9���9���9Į�9��9��9Ĵ�9k��9��9���9w��9���9̲�9���9԰�9���9¶�9��9��9���9#��9W��9���9���9x   x   ���9��9̯�9���9��9^��9a��9���9ϯ�9���9$��9Я�9\��9j��9ϳ�9o��9��96��9���9Ѱ�9ک�9��9ѭ�9è�9���9��9Գ�9���9��9���9x   x   ���9���9���9���9h��9?��9��9���9��9���9���9���9���9���9���9"��9���9`��9F��9���9��9���9ٳ�9���9̯�9��9m��9��9���9ʬ�9x   x   *��9k��9���9��9*��9��9���9���9հ�9���9h��9S��9��9ر�9��9���9c��9���9���9���9֭�9��9H��9���9���9��9 ��9a��9/��9;��9x   x   3��9۱�9ů�9س�9g��9|��9|��9��9J��9��9Ű�9[��9���9��9԰�9֬�9c��9���9T��9~��9Ĩ�9���9���9#��9z��9���94��9P��9@��9l��9x   x   .��9��9J��9;��9��9���9y��9P��9��9���9)��9
��9b��9���93��9���9n��9��9ʲ�9��9���9̯�9���9w��9���9ڲ�9X��9I��9���9J��9x   x   /��9���9���9|��9F��9̮�9���9���9��9ϰ�9��9���9;��9>��9}��9|��9���9"��9��9���9��9��9���9���9ز�9@��9۱�9_��9���9'��9x   x   ���9���9��9���9���9A��9���9@��9&��9Ѳ�9^��9W��9���9���9]��9���9J��9��9
��9#��9ӳ�9j��9���93��9X��9߱�9��9���9��9 ��9x   x   -��9Ѳ�9M��9{��9��9���9O��91��9į�9԰�9���9��9)��9���9���9Z��9s��9��9"��9V��9���9��9a��9N��9L��9b��9���9��9��9���9x   x   A��9m��9}��9���9ϳ�9N��9m��9��9ۭ�9��9B��9c��9���9���95��9l��9֮�9g��9L��9���9��9���92��9=��9���9���9��9��9
��9��9x   x   ۱�9���93��9%��9I��90��9���9��9x��9���9J��9��9,��9ï�9T��9֮�9a��9���9ڮ�9��9���9ʬ�9<��9o��9L��9'��9 ��9���9��9���9x   x   ���9r��9��9N��9ٷ�9��9��9y��9��9X��9���9;��9>��9���9δ�9��9��9���9U��9ı�9[��9��95��9\��9��9���9���9��9���9U��9x   x   y��9E��99��9m��9���9���9��9u��9���9���9��9���9Z��9g��9���9���9���9���9q��9��9���9��9B��9��9���9*��9е�9u��9M��9ݶ�9x   x   ��98��9���9.��9��9���9���9���9��9E��9��9��9u��9]��9��9���9��9��9���9���9���98��9��9[��9���9���9���9��9���9��9x   x   K��9l��91��9K��9���9���9϶�9���9��9���9U��9��9f��9���9���9A��9���9���9��9��9γ�9Ҷ�9y��9[��9{��9M��98��9��98��9۵�9x   x   ַ�9���9��9���96��9j��9���9p��9���9���9N��9	��9���9T��9j��9ɷ�9���9���9��9b��9���9@��9���9(��90��9ε�9���9ٷ�9��9��9x   x   ��9���9���9���9f��9ɲ�9Ե�9��9��9���9��9��9g��9¸�9���9���9��9��9���9���9��9E��9غ�9���9K��9��9��93��9��9E��9x   x   ��9��9���9Ӷ�9���9ص�9���9Ͷ�9���9&��9���97��9���9t��9ж�9��9(��9���9F��9��9���9C��9��9��9`��9���9V��9M��9l��9 ��9x   x   y��9x��9���9���9o��9��9Ͷ�9	��9'��9��9���9I��9���9߶�9ܺ�9=��9��9��9R��9���9m��97��9��9n��9���9��9���9̶�9��9���9x   x   ��9���9��9��9���9��9���9)��9��9��9S��9���9���9��92��9��9��9F��9F��9��9��9��9��9ĸ�9w��9���9H��9b��9:��9R��9x   x   V��9���9G��9���9���9���9%��9��9��9���9ӷ�9��93��9��9��99��90��9���9��9���9���9õ�9���9"��9B��9[��9��9&��9߷�9j��9x   x   ���9��9��9U��9M��9��9���9���9T��9ַ�9���9׷�9��9}��9Ե�9l��9���9��9���9���9��9��9��9��9���9s��9۶�9~��9R��9���9x   x   9��9���9��9��9
��9��96��9J��9���9��9۷�9���9Ķ�9���9���9T��9#��9��9F��9���9N��9
��9F��9���9��9��9϶�9���9%��9C��9x   x   =��9\��9p��9f��9���9d��9���9���9���95��9��9Ƕ�9ٴ�9N��9I��9õ�9c��9P��9��9д�9���9���9���9l��9���9���9��9r��9���9���9x   x   ���9i��9\��9���9Y��9���9v��9ݶ�9��9��9z��9���9Q��9��9c��9��9s��9���9X��9ٶ�9���9+��9���9��9D��9A��9��9��9���9���9x   x   ̴�9���9��9���9m��9���9ζ�9غ�9.��9��9ֵ�9���9I��9f��9U��95��9��9z��9з�9B��9���9s��9M��9���9��9I��9ϵ�9A��9���9���9x   x   ��9���9���9>��9Ʒ�9���9��9=��9��9:��9l��9R��9���9��96��97��9k��9d��9m��9Ͷ�9���9���9���9r��9Q��9��9���9���9��9��9x   x   ��9���9��9���9���9|��9'��9��9
��9,��9���9"��9f��9r��9��9k��9t��9���9۷�9��9���9���9i��9{��9��9X��9Ϸ�9���9��9��9x   x   ���9���9��9���9���9��9���9߶�9?��9���9��9��9V��9���9}��9d��9���9���9
��9��9���9��97��9���9ն�94��9{��9,��9���9,��9x   x   V��9u��9���9��9 ��9���9E��9R��9I��9	��9���9E��9
��9W��9ѷ�9i��9ڷ�9��9W��91��9���92��9��9¶�9��9(��9���9ָ�9d��9U��9x   x   ���9��9���9��9g��9���9��9���9��9���9���9���9ϴ�9׶�9C��9Ͷ�9��9��94��9��9>��9���9���9#��9v��9���9'��94��9k��9l��9x   x   [��9���9���9ϳ�9���9��9���9q��9��9���9��9O��9���9���9���9���9���9���9���9>��9���9F��9ʶ�9c��9���9ƴ�9Ŵ�9���9~��9"��9x   x   ��9��99��9Ѷ�9<��9C��9@��95��9��9ȵ�9��9��9���9+��9x��9���9���9��97��9ĸ�9K��9D��9س�9E��9��9ĵ�9q��9���9��9ڷ�9x   x   4��9B��9��9}��9Ż�9ߺ�9��9��9��9���9��9K��9���9���9P��9���9h��95��9��9���9ȶ�9ֳ�91��9E��9_��9!��9���9n��95��9��9x   x   _��9��9Z��9Z��9*��9���9��9s��9���9!��9߱�9���9k��9
��9���9m��9}��9���9���9��9]��9E��9G��9˸�9��9q��9���9���9ط�9���9x   x   |��9���9���9w��9-��9E��9\��9���9v��9B��9���9��9���9A��9��9V��9��9׶�9��9}��9���9��9]��9��9@��9���9
��9���9u��9Q��9x   x   ���9-��9���9L��9ѵ�9��9���9��9���9`��9p��9��9���9?��9M��9��9[��90��9'��9���9Ǵ�9µ�9!��9r��9���9o��9��9���9۴�9T��9x   x   ���9ѵ�9���98��9���9��9U��9���9I��9��9ض�9׶�9��9��9ε�9���9η�9}��9���9&��9Ĵ�9r��9���9���9	��9��9q��9<��9!��9y��9x   x   ��9u��9��9��9׷�94��9M��9϶�9a��9&��9~��9���9t��9��9A��9���9���9*��9ָ�93��9���9���9k��9���9���9���9>��9���9���9���9x   x   ���9K��9���93��9��9��9h��9��95��9߷�9Q��9'��9���9���9���9��9��9���9c��9l��9��9}��92��9ط�9s��9ٴ�9 ��9���9U��9���9x   x   X��9ݶ�9��9ص�9��9D��9"��9���9R��9h��9���9F��9���9���9���9��9��9+��9S��9n��9"��9ڷ�9��9���9S��9V��9z��9���9���9޶�9x   x   ��9��9���9���9d��9`��9x��9��9i��9I��9���9߿�9��9���9Ļ�9$��9���9o��9��90��9y��9Ⱦ�9"��9���9���93��9	��9��9��9���9x   x   ��9j��9y��9���9L��9���9���9���9��9ؽ�9x��9G��9۽�9���9���9���9u��9-��9���92��9��9��9f��9��9[��9��9���9��9��9���9x   x   ���9v��9`��9��9���9���9���9���9%��9���9޿�9&��9ػ�9h��9c��9/��9N��9Ի�9���9��9��9\��9���9���9���9���9���9��9���9��9x   x   ���9���9��9���9׽�9O��9��9���9y��9��9.��9��9j��9��9O��9���9���9���9��9м�9��9��9���9 ��9$��9X��9���9���9���93��9x   x   d��9J��9���9ս�9���9ѽ�9"��9{��9���9���9���9k��9½�9���9v��9E��9½�9��9��9���9���9#��9ӽ�9E��9��9��9��9Ѽ�9ؽ�9X��9x   x   ^��9���9���9S��9н�9���9M��9���9[��9н�9���9<��9۾�9��9w��9��9A��9��9���9��9���9Ƚ�9���9��9Q��9��9���9/��9��9Ͼ�9x   x   {��9���9���9���9!��9J��9��91��9p��9׽�9��9Y��9��9��9Ǿ�9��90��9<��9a��9���9���9\��9ѽ�9���9@��9���9��9w��94��9��9x   x   ��9���9���9���9{��9���92��9���9Ƚ�9Q��9���9���9���9(��9/��9���9u��9��9R��9���9��9���9���9���9��9˾�9 ��9���9���9ǿ�9x   x   j��9��9'��9|��9���9Y��9m��9ʽ�9���9���9��9^��9���9���9��9Խ�9��9��9���93��9k��9 ��9���9��9ʾ�9ƽ�9���9)��9��9g��9x   x   E��9Խ�9���9��9���9Ͻ�9Խ�9R��9���9���9Y��9ʽ�9���9���9!��9��9��9��9��9)��9���9���9���9���9��9���9u��9��9z��9��9x   x   ���9x��9޿�90��9���9���9��9���9��9W��9��9N��9=��9���9+��9��9���93��9���9���9���9���9C��9f��9d��9���9���9��9���9ƽ�9x   x   ��9E��9%��9��9h��9=��9[��9���9X��9Ž�9I��9P��9���9U��9	��9��9_��9Q��9q��94��9��9z��9!��9Z��9���9��9���9G��9	��9��9x   x   ~��9ܽ�9ۻ�9l��9½�9ܾ�9��9���9���9���9;��9���9���9���9R��9J��9P��9ڽ�9���9���9���9ۼ�9���9D��9���9N��9���9���9E��9U��9x   x   ���9���9g��9��9��9��9��9+��9���9���9þ�9R��9���9G��9C��9���94��9b��9ʿ�9���9���9��9ݾ�9��9ѿ�9r��9��9���9���9��9x   x   ���9���9e��9M��9x��9w��9ƾ�90��9��9 ��9*��9��9S��9D��9��9ӿ�9��9K��9˼�9P��9��9��9���9���9a��9���9u��97��9%��9��9x   x   "��9���9.��9���9C��9��9��9���9ս�9��9��9��9J��9���9ֿ�9N��9T��9��9��9���9���9x��9���9���94��9���9A��93��9v��9��9x   x   ���9r��9O��9���9½�9C��93��9r��9��9��9���9a��9M��9/��9��9R��9���9W��9��9���9e��9ݼ�9��9��9���95��97��9���9���9���9x   x   i��9,��9ѻ�9���9��9��9?��9��9��9��94��9P��9ٽ�9^��9J��9��9W��91��9s��9��9���9��9M��9���9_��9c��9��9���9A��9̻�9x   x   ��9���9���9��9��9���9f��9Q��9��9��9���9n��9���9ǿ�9ͼ�9��9 ��9x��9���9Ծ�9���9h��9���9��9���9���9���9м�9���9���9x   x   4��96��9��9Ҽ�9���9��9���9���92��9,��9���97��9���9���9Q��9���9���9��9Ӿ�9=��9D��9a��9ѻ�9Ⱦ�9l��9���9>��9&��9���9
��9x   x   |��9��9��9��9���9���9���9��9h��9���9���9��9���9���9��9���9`��9���9���9A��9F��9*��9��9���9���9���9Z��9���9>��9:��9x   x   ľ�9��9[��9��9%��9Ƚ�9^��9���9 ��9���9���9w��9ۼ�9��9��9v��9��9��9c��9^��9(��9ͽ�9���9ͼ�9���9_��9���9��9 ��9���9x   x   !��9g��9���9���9н�9���9ҽ�9���9���9���9E��9��9���9۾�9���9���9��9L��9���9һ�9 ��9���9���9���9c��9���9���9��9V��9���9x   x   ���9��9���9 ��9H��9��9���9���9��9���9g��9W��9G��9��9���9���9��9���9��9̾�9���9̼�9���9���9���9���9��9��9��9���9x   x   ���9Z��9���9#��9��9R��9>��9��9˾�9��9e��9���9���9տ�9c��9.��9���9a��9���9i��9���9���9f��9���9P��9x��9���9½�9���9,��9x   x   3��9��9���9W��9��9��9���9ʾ�9ƽ�9���9���9��9M��9p��9���9���9,��9g��9���9���9���9[��9���9���9y��9w��9���9Ѽ�9|��9���9x   x   ��9���9���9���9��9���9��9���9���9s��9���9|��9���9 ��9v��9F��98��9��9���9A��9]��9���9���9��9���9���9��9���9w��9���9x   x   ��9��9߽�9���9м�92��9w��9���9+��9��9��9B��9 ��9���95��97��9���9���9Ҽ�9&��9���9��9��9���9ý�9Ӽ�9���9���97��9��9x   x   ��9��9���9���9ܽ�9��93��9���9��9}��9���9��9G��9���9'��9z��9���9D��9���9���9<��9��9U��9��9���9~��9w��95��9ּ�9>��9x   x   ���9���9��95��9V��9Ҿ�9��9ǿ�9e��9��9ƽ�9��9U��9��9��9��9���9̻�9���9	��9:��9���9���9���9*��9���9���9��9=��9ƽ�9x   x   ���9
��9>��9��9}��9��9���9L��9��9���9���9���9D��9���9O��9���9-��9'��9���9���9���9���9���9���9���9���9��9���9$��9���9x   x   ��9���9���9@��9���9���9���9J��9���9'��9��9���9���9���9>��9��9���9���9���9���9���9k��9���9���9���9���9#��9l��9���9���9x   x   A��9���9���9���9 ��9���9���9Q��9���9���9���98��9F��9���9���9���9���9}��9���9���9���9m��9��9!��9���9&��9t��9��9���9���9x   x   ��9>��9���9|��9���9���9���9Q��9���9n��9���9���9���9z��9���9��9���9 ��9���9U��9|��9���9���9q��9���9'��9\��9���9���9\��9x   x   ��9���9 ��9���9���91��9���94��9d��9j��9���9���9���9B��9���9��9g��9"��9���9���9`��9���9���9���9���9���9\��9a��9���9���9x   x   ��9���9���9���90��9���9���9o��9��9���9���9��9���9���9���9���9���9 ��9 ��9���9e��9J��9���9��9���9��9��9���9	��9���9x   x   ���9���9���9���9���9���9��9���9`��9_��9���9��91��9A��9���9���9s��9*��9 ��9c��94��9���9e��9���9q��9��9���9���9���9���9x   x   L��9K��9Q��9T��96��9q��9���9N��9B��9]��9���9���9���9<��9��9��9���9d��9��9���9��9_��9 ��9���9{��9���9���9[��9��9���9x   x   ��9���9���9���9d��9��9b��9C��9���9���9 ��9���9\��9���93��9���9���9���9}��9���95��9��9��9���9���9)��9��9p��9���9���9x   x   ���9(��9���9l��9i��9���9^��9]��9���9G��9���9��9���9���9���9r��9S��9���9��9���9X��9���9���9Q��9U��9���9X��9���9���9l��9x   x   ���9��9���9���9���9���9���9���9%��9���9��9���9d��9T��9,��9>��9���9��9[��9���9���9}��9���9���9���9��9���9L��9���9���9x   x   ���9���99��9���9���9��9���9���9���9#��9���9p��9,��9A��9���9���9]��9���9���9���9���9���9;��9���9+��9��9I��9���9\��9��9x   x   H��9���9D��9���9���9���94��9���9a��9���9g��9*��9N��94��9}��9���9���9���9���9���9��9���9E��9g��9*��9���9���9���9g��9���9x   x   ���9���9���9~��9A��9���9>��9?��9���9���9W��9C��96��96��9���9���9���9Q��9��9a��9��9m��9%��9��9���9`��9���9���9���9���9x   x   O��9?��9���9���9���9���9���9��90��9���9,��9���9}��9���9%��9���9���9���9N��9_��9���9W��9���9>��9���9���91��9���9���9���9x   x   ���9��9���9!��9��9���9���9��9���9o��9?��9���9���9���9���9���9E��9��9��9c��9���9N��9���9���9���9X��9���9���9:��9R��9x   x   /��9���9���9���9c��9���9s��9���9���9Q��9���9Z��9���9���9���9D��9$��9���9���9"��9J��9p��9���9d��9���9���9���9��9���9��9x   x   +��9���9|��9���9 ��9��9'��9`��9���9���9��9���9���9X��9���9��9���9T��9���9T��9���9���9��9���9V��9���9��9���9���9���9x   x   ���9���9���9���9���9"��9��9��9~��9���9^��9���9���9��9J��9��9���9���9���9C��9���9���9/��9���9���9G��9���9p��9��9���9x   x   ���9���9���9X��9���9���9h��9��9���9���9���9���9���9]��9\��9d��9��9U��9C��9+��9���9��9w��9���9o��9���9���9%��9���9���9x   x   ���9���9���9~��9`��9a��97��9��96��9S��9���9���9~��9��9���9���9L��9���9���9���9���9���99��9^��9��9O��9���9���9)��9���9x   x   ���9n��9m��9���9���9L��9���9^��9��9���9���9���9���9p��9U��9O��9m��9���9���9���9���9���9t��9{��9_��9���9w��9>��9���9���9x   x   ���9���9��9���9���9���9e��9��9��9���9���9:��9I��9'��9���9���9���9��91��9y��97��9x��9���9��9X��9���9v��9p��9���9���9x   x   ���9���9#��9r��9���9��9���9���9���9O��9���9���9g��9��98��9���9b��9���9���9���9\��9{��9��9I��9���9c��9��9��91��9���9x   x   ���9���9���9���9���9���9t��9x��9���9R��9���9'��9*��9���9���9���9���9W��9���9o��9��9`��9W��9���9���9���9z��9���9��9/��9x   x   ���9���9%��9)��9���9��9��9���9-��9���9	��9��9���9c��9���9`��9���9���9J��9���9R��9���9���9d��9���9@��9���9N��9���9���9x   x   ��9"��9r��9]��9]��9��9���9���9��9X��9���9J��9���9���90��9���9���9��9���9���9���9v��9w��9��9{��9���9J��9���9t��9��9x   x   ���9q��9��9���9g��9���9���9Z��9o��9���9L��9���9���9���9���9���9��9���9l��9#��9���9<��9u��9��9���9I��9���9x��9���9���9x   x   "��9���9���9���9���9��9���9��9���9���9���9\��9g��9���9���99��9���9���9��9���9,��9���9���93��9��9���9t��9���9���9���9x   x   ���9���9���9\��9���9���9���9���9���9l��9���9"��9���9���9���9Q��9��9���9���9���9���9���9���9���92��9���9��9���9���9A��9x   x   R��9L��9��9���9���9���9	��9��9���9���9/��9���9���9��9<��94��9���9O��9/��9���9���9��9]��9���9���9���9���9���9���9I��9x   x   G��9��9n��9���9g��9Y��9���90��9���9x��9���9 ��9���9t��9��9F��9p��9���9���9���9���9���9^��9e��9���9M��9e��9��9��9���9x   x   ��9m��9R��9���9��9���9x��9���9���9W��9��9���9\��9���9���9��9���9���9���9���9���9Y��9���9��9���9���9���9���9��9]��9x   x   ���9���9���9���9���9���9���9���9
��9x��9���9K��9��9���9���9��9:��9���9���9`��9+��9���9���9���9���9;��9N��9���9��9��9x   x   ���9h��9 ��9���9U��9O��9?��9���9A��9���9��9���97��9m��9���9���9��9p��9��9���9���9 ��9y��9$��9P��9?��9���9��9���9G��9x   x   ���9[��9���9���9Q��9O��9f��9���9y��9E��9L��9]��9���9m��9���9���9z��9��9���9���9���9+��9��9.��9���9���9���9R��9���9���9x   x   ��9���9w��9���9B��9j��9d��9"��9R��9O��9���9���9���9
��9���9���9t��9���9_��9���9{��9!��9��9��9���9f��9���9���90��9+��9x   x   ��90��9���9���9���9���9��9S��9���9���9���9��9���9���9,��9��9���9���97��9(��9_��9o��9���9���9���9���9���9���9��9T��9x   x   ���9���9���9��9@��9y��9S��9���9���9���9��9���9��9���9���9R��9(��9��9���9���9���9���9���9���9b��9`��9���9���9���9��9x   x   ���9y��9Z��9{��9���9D��9O��9���9���9���9_��9���92��9���9���9}��9k��9���9��9X��9y��9���9���9���9���9���9c��9m��9���9J��9x   x   /��9���9��9���9��9J��9���9���9��9Y��9p��9C��9���9���9���9S��9��9D��9T��9=��94��9���9���9���97��9���9G��9��9R��98��9x   x   ���9��9���9L��9���9b��9���9��9���9���9@��9��9*��9���9��9?��9��9���9���9`��9 ��9���9���9~��9���9���99��9\��9#��9���9x   x   ���9���9\��9��92��9���9���9���9��92��9���9'��9n��9S��9��9���9���9��94��9���9���9k��9���9��9M��9���9���9���9���9\��9x   x   ��9u��9���9���9j��9l��9	��9���9���9���9���9���9X��9'��9���9���9G��9���9���9���9���9���9 ��9Q��9J��9���9���9��9V��9��9x   x   A��9��9���9���9���9���9���90��9���9���9���9��9��9���9w��9���9���9g��9 ��9_��94��9o��9���9l��9.��9���9)��9���9��9���9x   x   7��9G��9��9��9���9���9���9��9U��9���9V��9=��9���9���9���9���9���9��9=��9X��9r��9r��9y��9��9���9���91��9V��9���99��9x   x   ���9n��9���9:��9��9y��9w��9���9'��9j��9��9��9���9C��9���9���9���9���9S��9���9���9��9p��9��9r��9���9���9���9���9��9x   x   M��9���9���9���9t��9��9���9���9��9���9G��9���9��9���9e��9���9���9���9���9���9:��9��9��95��9���9���9���9%��9t��96��9x   x   -��9���9���9���9��9���9\��94��9���9��9U��9���92��9���9#��9=��9T��9���9_��9���9���9*��9���9���9���9F��9��9���9���9���9x   x   ���9���9���9^��9���9���9���9(��9���9S��9<��9`��9���9���9b��9W��9���9���9���9#��9���9���9���9���9���9y��9���9���9Y��9���9x   x   ���9���9���9*��9���9���9v��9_��9���9{��95��9��9���9���92��9r��9���9:��9���9���9���9Y��9L��9��9���9���9'��9���9-��96��9x   x    ��9���9W��9���9 ��9'��9!��9l��9���9���9���9���9j��9���9l��9p��9	��9��9"��9���9\��9��9���9o��9���9+��9���9���93��9���9x   x   ]��9_��9���9���9|��9��9	��9���9���9���9���9���9���9���9���9x��9r��9��9���9���9K��9���9���9G��9���9���9���9���9=��9���9x   x   ���9e��9��9���9$��90��9��9���9���9���9���9}��9��9T��9n��9��9��9/��9���9���9��9q��9F��9���9���9���9���9���9���9T��9x   x   ���9���9���9���9M��9���9���9���9e��9���98��9���9P��9L��9.��9���9s��9���9���9���9���9���9���9���9��9���9���9��9q��9��9x   x   ���9P��9���9=��9C��9���9g��9���9a��9���9���9���9���9���9���9���9���9���9D��9w��9���9,��9���9���9���9���9���9W��9���9���9x   x   ���9c��9���9K��9���9���9���9���9���9c��9F��9;��9���9���9%��9.��9���9���9��9���9$��9���9���9���9���9���9���9��9/��96��9x   x   ���9��9���9���9��9V��9���9���9��9m��9��9^��9���9��9���9Z��9���9(��9��9���9���9���9���9���9��9Y��9 ��9P��9���9%��9x   x   ���9��9��9��9���9���92��9��9���9���9M��9"��9���9W��9��9���9���9u��9���9W��9.��92��9<��9���9r��9���9/��9���9Z��9���9x   x   I��9���9]��9��9I��9���9.��9S��9��9K��98��9���9Z��9��9���9<��9��9<��9���9���97��9���9���9R��9��9���95��9&��9���9W��9x   x   c��9���9��9���9��9Q��9n��9���9 ��9U��9���9?��9���9(��9���9���9��9���9��9\��9���9���9���9���9���9���91��9���9���9���9x   x   ���9���9���94��9���9��9���9��9r��95��9���9��9��9v��9!��9���9Y��9e��9J��9���9���95��9%��9���9���9���9'��9��9���9���9x   x   ���9���9��9���9{��9r��9���9���9 ��9e��9J��9x��9g��9���9��9���9���9���9���9��9r��9T��9y��9���9���9��9_��9Y��9��9j��9x   x   ���96��9���9w��9"��9���9C��9L��9,��9��9���9���9l��9~��9���9���94��9���9���9���9���9���9���93��9~��9���9I��9J��9t��9/��9x   x   
��9���9x��9#��9���9��9/��9/��9���9���9n��9���9���9���97��9���9z��9��9Q��9���9��9f��9M��9e��9��9d��9B��9���9���9���9x   x   N��9��9r��9���9��9���9u��9���9i��94��9���9���9h��9$��9���9*��9���9;��9���9)��9��9���9 ��9h��9=��9K��9���9���9���9g��9x   x   q��9���9���9A��9,��9s��9��9#��94��9���9���9��9H��9|��9���9���9���9��9���9}��9r��9d��9#��9$��9I��9���9��9E��9���9��9x   x   ���9��9���9K��9/��9���9!��9���9���9R��9n��9��9��9P��9|��9P��9��9'��9��99��9R��9���9��9?��9���9���9i��9���9���9=��9x   x   &��9t��9��90��9���9j��95��9���9���9
��9z��9m��9���9��9���9���9(��9���9Q��9��9S��9���9��9)��9���9���9��9R��9���9���9x   x   U��92��9d��9��9���94��9���9T��9
��9Z��9P��9!��9��9���9���9��9z��9.��9���9	��9��9e��9g��9���9���9Q��9���9>��9���9��9x   x   ���9���9F��9���9n��9���9���9n��9|��9V��9V��9H��9���9��9���9\��9���9[��9���9w��9C��9���9���9y��9���99��9���9g��9P��9Q��9x   x   E��9��9y��9���9���9���9��9��9p��9(��9F��9���9���9��9���9���9-��9���9W��9���9(��9���9m��9���9s��9Z��9��9���9���9���9x   x   ���9��9l��9j��9���9h��9I��9��9���9��9���9���9���9���9z��9��9T��9���9��9���9���9���9��9���9���9���9���9���9���9U��9x   x   *��9r��9���9~��9���9#��9~��9Q��9��9���9��9��9���9 ��9���9t��9���9���9���9���9e��9W��9^��9���9���9���9'��9<��9���9��9x   x   ���9��9��9���9:��9���9���9z��9���9���9���9���9{��9���9g��9	��9a��9<��9O��9���9���95��9���9��9���9l��9���9��9���9E��9x   x   ���9���9���9���9���9(��9���9H��9���9��9[��9���9��9s��9��9���9���9���9���9��92��9���9���9���9��9i��9���9���9���9���9x   x   ��9X��9���99��9x��9���9���9��9%��9w��9���90��9U��9���9e��9���9��9Z��9���9g��9��98��9���9W��9D��9���9@��94��9���9���9x   x   ���9h��9���9���9��99��9��9(��9���9.��9Z��9���9���9���9:��9���9X��9���9���9���9���9���9#��9��9~��9P��9���9^��9`��9=��9x   x   ��9L��9���9���9T��9���9���9��9R��9���9���9U��9��9���9N��9���9���9���9���9;��9(��9g��9���9��9���9���9���9���9-��9��9x   x   ^��9���9��9���9���9(��9~��97��9��9��9y��9���9���9���9���9��9h��9���9<��9?��9���9���9���9]��9���9"��9��9���9���9���9x   x   ���9���9s��9���9��9��9u��9V��9Q��9��9A��9%��9���9g��9���9/��9��9���9*��9���9*��9I��9���9���94��9!��9*��9o��9���9p��9x   x   ���92��9S��9���9h��9���9e��9���9���9d��9���9���9���9Y��99��9���9;��9���9g��9���9J��9���9��90��9D��9���9���9"��9P��9���9x   x   ���9$��9|��9���9I��9���9!��9��9��9i��9���9o��9��9^��9���9���9���9%��9���9���9 ��9��9���9��9B��9���9���9��9
��9A��9x   x   ���9���9���96��9f��9h��9#��9?��9&��9���9u��9���9���9���9��9���9W��9$��9��9^��9���9.��9��9���9���9��9���9���9��9���9x   x   ���9���9���9���9��9;��9G��9���9���9���9���9u��9���9���9���9��9F��9}��9���9���97��9C��9D��9���9��9���9���9���9n��9:��9x   x   ���9���9��9���9f��9M��9���9���9���9R��99��9Y��9���9���9m��9h��9���9P��9���9��9#��9���9���9��9���9.��9g��9���9���9���9x   x   0��9*��9b��9H��9E��9���9��9l��9��9���9���9��9���9,��9��9���9A��9���9���9��9,��9���9���9���9���9e��9���9���9��9���9x   x   ���9��9\��9G��9���9���9C��9���9O��9?��9i��9���9���99��9��9���91��9\��9���9���9m��9"��9��9���9���9���9���9���9���9��9x   x   ���9���9��9u��9���9���9���9���9���9���9O��9���9���9���9���9���9���9_��9*��9���9���9S��9��9��9n��9���9���9���9L��9���9x   x   ���9���9i��90��9���9f��9��9;��9���9��9T��9���9Y��9��9D��9���9���9<��9��9���9n��9��9?��9���9;��9���9���9}��9���9���9x   x   ���9&��9��9 ��9T��9;��9���92��9���9���9���9{��9���9���9Q��9��9���9T��9���9`��9Y��9g��9��9@��9���9��9��9 ��9���9O��9x   x   $��9���9��9P��9���9?��9 ��9���9N��9���9P��9���9���9���9���9���9���9���9���9���9��9
��9e��9���9���9���9���9���9z��9E��9x   x   ��9��9M��9��9��9���9{��9���9U��9���9��9���9i��9���9z��9���9���9/��9���9X��9���9��9���9+��9���9g��9���9V��9��91��9x   x   ��9N��9��9R��9���9���9��9���9��9'��9\��9���9:��9h��90��9���9���9���9��9���93��9���95��9���9��9
��9
��9���9/��9���9x   x   U��9���9��9���9��9(��9J��9���9x��9q��9���9���9���9w��9@��91��9 ��9=��9m��9f��9���9��9o��9���9
��9Y��9^��9���9���9��9x   x   =��9>��9���9��9&��9l��9��9d��9 ��9{��9���9���9���9���9���94��9=��9Q��9���9���9{��9���9���9 ��9��9C��9d��9���9r��9���9x   x   ���9��9}��9��9L��9��9��9���9���9X��9���9e��9���9T��9���9��9���9+��9p��9���9���9n��9X��9?��9���9h��9y��9���9*��9R��9x   x   0��9���9���9���9���9e��9���9T��9���9:��9e��90��9���9n��9���9���9���9���9F��9���9���9Z��95��9���9���9���9\��9���9���9���9x   x   ���9N��9S��9��9v��9!��9���9���9��9���9,��9���9_��9���9���9k��9���9���9^��9���9��9z��9I��9-��9��9���9���9���9���9%��9x   x   ���9���9���9%��9p��9y��9^��9:��9���9��9���9��9���9���9���9a��9\��9���9���9{��9?��9���9��90��9���9���9��9��9���9D��9x   x   ���9P��9��9^��9���9���9���9a��9+��9���9��9���9r��9���9��9���9���9-��9���9���9@��9W��9���9O��9i��9#��9���9���9���9���9x   x   y��9 ��9���9���9���9���9f��9-��9���9��9���9'��9���9���9��9���9x��9���9v��9���9H��9���9A��9���9i��9@��9p��9��9!��9��9x   x   ���9���9i��99��9���9���9���9���9^��9���9r��9���9���9\��9K��9���9x��9���9��9��9���98��9F��9���98��9���9���9���9���9��9x   x   ���9���9���9g��9{��9���9R��9m��9���9���9���9���9W��9A��9���9���9���9X��9���9l��9.��9~��9���9���9y��9���9J��9���9���9w��9x   x   T��9���9{��9-��9A��9���9���9���9���9���9��9%��9K��9���9���9^��9i��9��9���9V��9���9���99��9o��9���9B��9���9���9���9���9x   x   ��9���9���9���91��94��9
��9���9u��9a��9���9���9���9���9^��9y��9��9���9W��9���9���9j��9z��9)��9M��9���9���9��9`��9���9x   x   ���9���9���9���9!��9?��9���9���9���9_��9���9{��9v��9���9d��9}��9���9��9L��9B��9���9y��9���9���9x��9��9���9���9@��9���9x   x   W��9���90��9���9=��9O��9)��9���9���9���9*��9���9���9Z��9��9���9��9���9���9c��9���9���9<��9���9���9��9���9?��9���9=��9x   x   ���9���9���9��9l��9���9q��9H��9^��9���9���9u��9|��9���9���9X��9H��9���9���9���9$��9���9}��98��9���9���9���9���9"��9D��9x   x   _��9���9Z��9���9h��9���9���9���9���9{��9���9���9��9i��9V��9���9A��9d��9���9���9��9��9���9���9���91��9���9���9[��9_��9x   x   W��9��9���95��9���9u��9���9���9
��9=��9>��9K��9���9,��9���9���9���9���9#��9��9b��9��9���9s��9���9���9��9���9��9���9x   x   k��9��9��9���9��9���9k��9\��9|��9���9Z��9���95��9|��9���9n��9z��9���9���9!��9��9���9O��9���9���9���9���9���9���9��9x   x   ��9h��9���95��9p��9 ��9W��97��9K��9��9���9A��9H��9���96��9|��9���95��9{��9���9���9M��9-��9a��9��9F��9l��9���9|��9���9x   x   @��9���9)��9���9���9"��9=��9���9/��9-��9N��9���9���9���9q��9*��9���9���98��9���9r��9���9c��9 ��9U��9���9U��9w��90��9���9x   x   ���9���9���9��9��9��9���9���9��9���9i��9e��97��9x��9���9N��9x��9���9���9���9���9���9��9T��9���9���9���9���9O��9R��9x   x   ��9���9e��9
��9Q��9A��9f��9���9���9���9"��9@��9���9���9A��9���9��9��9���92��9���9���9C��9���9���9���9��9h��9��9T��9x   x   	��9���9���9��9`��9g��9v��9b��9���9��9���9n��9���9G��9���9��9���9���9���9���9��9���9k��9S��9���9��9t��9���9���9���9x   x   !��9���9X��9���9���9���9���9���9���9��9���9��9���9���9���9��9���9=��9���9���9���9���9���9v��9���9g��9���9{��9z��9���9x   x   ���9x��9��9,��9���9r��9*��9���9���9���9���9��9���9���9���9f��9F��9���9'��9b��9��9���9~��92��9Q��9��9���9}��9^��9���9x   x   S��9I��92��9���9��9���9R��9���9(��9E��9���9��9��9x��9���9���9���9:��9E��9a��9���9��9���9���9S��9X��9���9���9���9C��9x   x   ��9���9��9���9O��9���9���9���9���9���9���9���9��9���9���9��9V��9���9���9���9���9���9m��9e��9m��9���9���9R��9���9���9x   x   ���9���9���9Q��9 ��9��9���9��9��9!��9X��9E��9<��9��9��9��9c��9k��9���9��9���9��9���9���96��95��9���9$��9���9q��9x   x   ��9���9���9���9 ��9���9o��9B��9���9���9D��9��9}��9R��9���9}��9���9���9t��9���9���9���9���9��9���9^��9���9U��9��9���9x   x   ���9O��9���9v��99��9w��9���9J��9���9���9���9"��9���9���9���9��9���9���9B��9���9���9+��9���97��9F��9���9���9a��9���9���9x   x   P��9���9��9:��9v��99��9p��9D��9"��9���9��9>��9��9���9���9��9���9���9���9X��9���9���9Y��9���9���9���9���9V��9=��9���9x   x   ���9���9���9v��9=��9g��9���9���9��9��9��9���9���9i��9I��9���9[��9���9&��97��9Y��9��9���9K��9|��9c��9e��9V��9���9���9x   x   ���9���9o��9���9p��9���9���9��9*��9���9)��9A��9���9{��9���9���9���9���9���9��9��9���9���9���9��9��9���9���9���9!��9x   x   ���9��9D��9I��9B��9���9��9���9o��9���97��9���9���9���9+��9���9n��9��9���9���9^��9���9���9&��9���9���9���9���9���9���9x   x   ���9��9~��9���9%��9��9+��9n��9���9G��9���9���9���9���9���9���9o��9I��9���9���9���9���9 ��9��9���9���9���9��9)��9R��9x   x   ���9$��9���9���9���9���9���9���9I��9���9��9���9���9���9s��9��9���9
��9T��9���9���9���9r��9n��9S��9���9G��9���9x��9���9x   x   ���9Y��9B��9���9��9��9-��98��9���9��9y��9��9���9$��9���9n��92��9���9F��9"��9���9���9���9���9���9t��9��9'��9��9���9x   x   ���9C��9��9"��9@��9���9F��9���9���9���9��9���9���9���9���9`��9{��9��9���9���9���9���9Y��99��9��9J��9[��9!��9���9���9x   x   ��9=��9}��9���9��9���9���9���9���9���9���9���9W��9L��9���9y��9^��9���9e��9���9A��9!��9��9��9/��9���9���9���9��9���9x   x   ���9��9N��9���9���9k��9}��9���9���9���9#��9���9L��9���94��9V��9���9F��9W��9���9���9)��9���9���9q��9���9���9S��9>��9/��9x   x   ���9��9���9���9���9F��9���9,��9���9t��9���9���9���97��9(��9m��9X��9q��9���9���9���9���9��9��9}��9���9���9���9���9"��9x   x   ��9��9~��9��9��9���9���9���9���9��9m��9_��9{��9Y��9n��9���9���9���9���9���9���9���9���9���9z��9A��9���9���9���9#��9x   x   W��9h��9���9���9���9[��9���9n��9i��9���95��9|��9`��9���9Y��9���9
��9��9���9��9���9^��9���9d��95��9���9���9���9��9���9x   x   ���9k��9���9���9���9���9���9��9I��9��9���9��9���9G��9o��9���9��9r��9���9��9���9	��9��9���9���9@��9���9^��9���9���9x   x   ���9���9r��9C��9���9$��9���9���9���9S��9G��9���9c��9Z��9���9���9���9���9���9���9���9d��9���9���9_��9K��90��9���9���9���9x   x   ���9��9���9���9X��99��9"��9���9���9���9"��9���9���9���9���9���9��9"��9���9���9}��9���9��9j��9���9���90��9���92��9���9x   x   ���9���9���9���9���9\��9��9a��9���9���9���9���9A��9���9���9���9���9���9���9u��9s��9���9���9���9��9���9���9~��9���9X��9x   x   ���9��9���9,��9���9��9���9���9���9���9���9���9#��9-��9���9���9\��9��9d��9���9���9
��9P��9}��9���9���9���9(��9���9S��9x   x   h��9���9���9���9X��9���9���9���9��9m��9���9\��9��9���9��9���9���9��9���9��9���9P��9^��9���9���9W��9P��9^��9{��9���9x   x   g��9���9���95��9���9J��9���9#��9��9k��9���99��9��9���9��9���9j��9���9���9m��9���9���9���9%��9���9���9���9>��9���9H��9x   x   k��97��9���9G��9���9���9��9���9���9V��9���9 ��9.��9p��9���9x��92��9���9`��9���9��9���9���9���9���9���9Y��9���9���9>��9x   x   ���99��9b��9���9���9c��9��9���9���9���9s��9N��9���9���9���9=��9���9@��9K��9���9���9���9Y��9���9���9��9��9R��9���9���9x   x   ���9���9���9���9���9e��9���9���9���9H��9��9X��9���9���9���9���9���9���92��9.��9���9���9Q��9���9W��9!��9��9��9<��9d��9x   x   R��9&��9R��9`��9U��9Y��9���9���9��9���9)��9$��9���9Z��9���9���9���9^��9���9���9���9'��9b��9;��9���9T��9��9��9��9���9x   x   ���9���9��9���9;��9���9���9���9-��9u��9��9���9 ��9<��9���9���9	��9���9���9-��9���9���9~��9���9���9���9:��9��9��90��9x   x   ���9p��9���9���9���9���9 ��9}��9Q��9���9���9���9���9-��9&��9"��9���9���9���9���9^��9R��9���9D��9;��9���9_��9���9.��9���9x   x   ��91�9��9%	�9�9��9��9u�9
�9��9�	�9e�9b�9�	�9��9^�9}�9
�9��9��9;	�9�9��9��9��9{�9�9��9��9J�9x   x   -�9t�9	�9��9��9��9�9&�9��9��9��98�9@�9A�9��9��9B�9��9��9�9��9/	�9i	�9��9�9{�9o�9��9��9'�9x   x   ��9	�9�
�9��9��9N�9,	�9}�9�9j�9�
�9��9o�9;�9��9M�9��9�9�
�9y�9��9q�9��9S�9��9l�91�9�	�9K�9�	�9x   x   !	�9��9��96�9�9	�9+�9��9��9�	�9�	�9��9��9x�9��9��9��9�	�9	�9`�9�	�9:�9�	�9��9��9��9J�9�	�9��9��9x   x   ~�9��9��9�9��9��9��9
�96	�9��9u�9��9	�9��9��9�9��9	�9�	�9�	�9��9��9��9/�9�9��9Z�9�9��9^�9x   x   ��9��9P�9	�9��9��9V	�9)	�9�9+�9��9	�9��9)�9��9��9�9��92	�95	�9:	�9��92	�9��94�9��9&�9#	�9��9�9x   x   ��9�9+	�9)�9��9[	�9;�9��9e�9`�9�9�	�9V�9�	�9
�97�9��9�9��9��9��9��9��9��9s�9��9��9��9�9��9x   x   r�9 �9��9��9
�9*	�9��9{�9��9v	�9��9��9��9%�9
�9O�9�9��90	�9�
�9�9��9�93�9�
�9�94	�9B	�9�
�9$
�9x   x   
�9��9�9��94	�9�9i�9��9Z
�9��9?�9
	�9��9	�9
�9X�9X�94�9n	�9>�9��9V	�9�	�9A�9�9�9��9�9y�9T�9x   x   ��9��9i�9�	�9��9/�9]�9u	�9��9N�9�
�9�
�9c�9�9�
�9��9�9�	�9I�9��9��9��9$	�9��9��9�	�9�	�9��9��9U�9x   x   �	�9��9�
�9�	�9u�9��9�9��9>�9�
�9��9�
�9��9��9z
�9�9��9R
�9�
�9��9
�9L	�9/�95�9��9��9��9�94�9	�9x   x   j�9:�9��9��9��9�9�	�9��9	�9�
�9�
�9I�9��9�	�9�9s�9��95�9��9�9;�9P�9��9w�9��9��9��9�96�9%�9x   x   `�9?�9n�9��9
�9��9N�9��9��9`�9��9��96�9Z�9�9t�9��9 �9�9��9�	�9�	�9��9��9��9H�9[�98
�9
�9�9x   x   �	�9A�9;�9{�9��9/�9�	�9 �9��9�9��9�	�9]�9^�9��9�9p�9�	�9�
�9��9r�9=	�9l�9�9�9�9��9d�9��9�
�9x   x   ��9��9��9��9��9��9
�9
�9
�9�
�9z
�9�9�9��9��9r�9��9 �9��9��9X�9_�9�9��9��9��9[�9��9��9�9x   x   _�9��9G�9��9 �9��9<�9T�9Y�9��9�9s�9t�9�9o�9k�9��9i	�9��9 	�9�	�9;�9�
�9�	�9N�9
�9��9]�9�	�9|�9x   x   ��9C�9��9��9��9�9��9�9W�9�9��9��9��9r�9��9��9��9.�9��91�9x�9Q
�9�
�9=�9�
�9��9�	�9�9$	�9j�9x   x   
�9��9�9�	�9	�9��9�9��96�9�	�9R
�92�9�9�	�9�9i	�90�9��9��9��9��9U�9}�9��9��9 �9��9��9�	�9'�9x   x   ��9��9�
�9	�9�	�93	�9��9/	�9s	�9L�9�
�9��9�9�
�9��9��9��9��9��9�	�9U�9��9��9
�9��9t�9�	�9b�9��9�
�9x   x   ��9�9u�9e�9�	�96	�9��9�
�9=�9��9��9�9��9��9��9 	�91�9��9�	�9��9B�9��9��9��9t	�9��9��9��9I	�9��9x   x   <	�9��9��9�	�9��9<	�9��9�9��9��9
�9<�9�	�9m�9X�9�	�9w�9��9Y�9D�9`
�9p�9��9Z�9Y�9�	�9��9��93
�9F�9x   x   �90	�9q�9:�9��9��9��9��9R	�9��9O	�9P�9�	�9@	�9b�9?�9N
�9Q�9��9��9p�9��9��9|
�9��9�9D	�9+
�9�9�	�9x   x   ��9l	�9��9�	�9��90	�9��9�9�	�9)	�94�9��9��9l�9�9�
�9�
�9z�9��9��9��9��9��9�	�9�9L�9��9��9	�9	�9x   x   ��9��9U�9��96�9��9��94�9?�9��93�9w�9��9�9��9�	�99�9��9
�9��9[�9y
�9�	�9*�9[�9�9C�9��9��9��9x   x   ��9�9��9��9�91�9t�9�
�9�9��9��9��9~�9�9��9P�9�
�9��9��9w	�9[�9��9�9\�9P�9��9P�9��9��9�
�9x   x   z�9{�9f�9��9��9��9��9�9�9�	�9��9��9I�9�9��9
�9��9�9t�9��9�	�9
�9M�9�9��9C�9k	�9��9U
�9H�9x   x   �9r�91�9L�9\�9%�9��95	�9��9�	�9��9��9\�9��9Y�9��9�	�9��9�	�9��9��9>	�9��9G�9T�9j	�9�9!	�9�9��9x   x   ��9��9�	�9�	�9�9	�9��9B	�9�9��9�9 �94
�9b�9��9^�9�9��9c�9��9��9+
�9��9��9��9��9	�9Y�9��9L�9x   x   ��9��9O�9��9��9��9�9�
�9y�9��94�97�9
�9��9��9�	�9%	�9�	�9��9J	�93
�9�9�9��9��9U
�9�9��9�	�9H�9x   x   F�9$�9�	�9��9^�9�9��9$
�9V�9X�9	�9)�9�9�
�9�9��9n�9+�9�
�9��9J�9�	�9��9��9�
�9E�9��9L�9D�9K	�9x   x   ��9;�9=�9�9��9��9s�9��9��9��9=�9�9��99�9��9i�9��9C�9��9��9��9��95�90�9)�9
�9��9@�9V�9E�9x   x   :�9��9��9��9[�9��9O�9!�9�9�9B�9R�9��9��9q�9�9s�9��9<�90�9h�9"�9B�9��9��9��9��9��9��9��9x   x   >�9��9T�9N�9%�9��9��99�9f�9�9��9C�9��9��9�9J�9��9V�9T�9,�9��95�9��9�9��9?�9��9u�9y�9��9x   x   �9��9Q�96�9q�9&�9�9��9��9n�9��9��9��9}�9h�9��9l�9!�9��9��9��9�9w�9{�9@�9�9��9��9%�9��9x   x   ��9Y�9#�9q�9N�9��9��9��9��9�9��9��9��97�9��9��9��9{�9��9��9��9��9��9��9p�9��9��9G�9��93�9x   x   ��9��9��9#�9��9&�9\�9+�9��9�9k�9	�9�9��9��9��9>�9��9K�9M�9|�9�9��9��9��9��9P�9��9;�9��9x   x   t�9Q�9��9�9��9[�97�9�9$�9��9��9��9�9��9��9��9�9U�9��9�9�9�9��9��9�9��9��9�9N�9��9x   x   ��9!�97�9��9��9,�9�9T�9��9��9 �9��9��9�98�9(�9��9��9��9��9��9��9\�9�9��9�96�9�9�9��9x   x   ��9�9c�9��9��9��9�9��9�9��9`�9��9�9�9��9#�9��9��9��92�9��9}�9��9�9�9l�9��9��9*�9��9x   x   ��9�9�9n�9�9�9��9��9��9�9��9��9[�9��9��9��91�9�9Y�9�9��9��9��9�9Q�9��9��9��9��9<�9x   x   ;�9A�9��9��9��9l�9��9�9^�9��9��9��96�9��9%�94�9��9��9��9�9R�9@�9��9:�9��9��9j�9�9��9��9x   x   �9P�9A�9��9��9�9��9��9��9��9��9��9��96�9�9^�9��9��9��9��9��9I�9v�9��9K�9�9*�9.�9�9��9x   x   ��9��9��9��9��9�9�9��9�9[�96�9��9 �9&�9w�9T�9G�9b�9�9�9��9��9��9��9��9��9��9u�9��9��9x   x   =�9��9��9y�97�9��9��9 �9��9��9��93�9#�9��9��9��9��9�9�9K�9F�9�9 �9��9=�9��9��9��9��9��9x   x   �9o�9��9h�9��9��9��94�9��9��9!�9�9x�9��9��9L�9m�9��9��9�9�9�9g�9��9��9��9��9��9s�9��9x   x   l�9�9P�9��9��9��9��9+�9"�9��93�9_�9W�9��9N�9��9��95�9t�9�9g�9]�9��9 �9N�9+�9��9��9��9m�9x   x   ��9o�9��9j�9�9=�9
�9��9��9/�9��9��9G�9��9j�9��9��9�9�9P�9m�9�9]�9��9R�9��9��9Q�9*�9D�9x   x   E�9��9X�9%�9w�9��9P�9��9��9	�9��9��9c�9�9��95�9�9��9G�9��9��9G�9y�9n�9��9��9��9��9��9��9x   x   ��9:�9X�9��9��9N�9��9��9��9X�9��9��9�9�9��9v�9��9G�9*�9��9#�9,�9d�9��9��9K�9��9:�97�9E�9x   x   ��93�9+�9��9��9O�9�9��91�9�9�9��9�9I�9�9�9P�9��9��9�9��9I�9�9%�9��9��9��9��9��9��9x   x   ��9i�9��9��9��9w�9�9��9 �9��9S�9��9��9G�9�9f�9m�9��9"�9��9��9)�9��9�9��98�9��9]�9��9�9x   x   ��9"�94�9�9��9#�9�9��9~�9��9=�9G�9��9�9�9[�9�9E�9*�9H�9'�9��9�94�9��9��93�96�9�9��9x   x   8�9A�9��9u�9��9��9��9Z�9��9��9��9u�9��9�9d�9��9a�9y�9f�9 �9��9�99�9~�9%�9�9�9��9��9��9x   x   /�9��9�9x�9��9��9��9�9�9�9;�9��9��9��9��9�9��9o�9��9(�9�94�9��9O�9�9b�9-�9�9��9��9x   x   +�9��9��9A�9s�9��9
�9��9�9S�9��9G�9��9>�9��9N�9Q�9��9��9��9��9��9&�9�9��9��9��9`�9'�9��9x   x   
�9��9@�9~�9��9��9��9�9h�9��9��9�9��9��9��9+�9��9��9M�9��9:�9��9�9c�9|�9
�91�9��9@�9��9x   x   ��9��9��9��9��9R�9��96�9��9��9l�9(�9��9��9��9��9��9��9��9��9��97�9	�90�9��9.�9��9x�9��9��9x   x   ?�9��9s�9��9I�9��9�9�9��9��9�9-�9x�9��9��9��9N�9��9:�9��9]�9=�9��9	�9b�9��9x�9��9��9�9x   x   V�9��9y�9$�9��9<�9L�9�9*�9��9��9�9��9��9x�9��9)�9��98�9��9��9�9��9��9%�9A�9��9��9��9��9x   x   J�9��9��9��95�9��9��9��9��9@�9��9��9��9��9��9h�9B�9��9B�9��9�9��9��9��9��9��9��9�9��9��9x   x   k1�9,�9�*�9�,�9n+�9�*�9�*�9+�9,�9�,�9�)�9�(�9�*�9�'�9�(�9�&�9�&�9�*�9�*�9q)�9�)�9w+�9�+�9s+�9+�9�)�9�,�9-�9�*�9,�9x   x   ,�9K.�9�,�9E,�9(�9�(�9-�9�+�9D-�9>+�9�)�9],�9a,�9)(�9�(�9�*�9'�9�*�9�+�9)�9�,�9�-�9,�9K,�9�(�9�'�9z+�9r,�9�.�9�,�9x   x   �*�9�,�9�)�9�(�9�*�9�(�9Y*�9�*�9*�9�+�9�,�9$*�9-�9�-�9�*�9�-�9m-�9�+�9m-�9�*�9l)�9T*�9�*�9 )�9!+�9�(�9y*�9:-�9*�9W%�9x   x   �,�9A,�9�(�9-,�9�,�9�)�9�-�9f*�9�,�9�,�9+�9^*�9�'�9�'�9�%�9�(�9n)�9)�9�-�9-�9.+�9�-�9�)�9�+�9�,�9�(�9�*�9/-�9/�9�.�9x   x   o+�9(�9�*�9�,�9�+�9�+�9�,�9�,�9.�9:)�9)+�90+�9o*�9�,�9�+�9S*�9A-�9P)�9B-�9k,�9�,�9�+�9J,�9�,�9J*�9G)�9,�9+�9G,�9/,�9x   x   �*�9�(�9�(�9�)�9�+�9U(�9�*�9O+�9�+�9�+�9�'�9,�9�,�9�,�9+�9�'�9�*�9�+�9],�9�*�9t(�9�*�9J)�9)�9�(�9~)�9i-�9'(�9]'�9-�9x   x   �*�9-�9[*�9�-�9�,�9�*�9&(�9�(�9�*�9�)�9�*�9�,�9q(�9�,�9�,�9I(�92,�9(�9�'�9�*�9�,�9.�9*�9�,�9F+�9(,�93-�9b-�9�-�9Q+�9x   x   +�9�+�9�*�9i*�9�,�9N+�9�(�9�/�9�+�9 *�9�/�9�)�9*�9K.�9=*�9o,�9�.�9t)�98+�9�,�9�)�9�*�9�+�9�*�9�(�9�'�9�)�9�)�9�(�9')�9x   x    ,�9A-�9*�9�,�9.�9�+�9�*�9�+�9�&�9�+�9�-�9T&�9�.�9�+�9�&�94+�9�+�9�+�9+.�9U-�9�)�9P-�9S,�9�+�9�*�9�,�9-�9z+�9*�9�+�9x   x   �,�9F+�9�+�9�,�99)�9�+�9�)�9*�9�+�9Y/�9Y+�9�)�9�/�9,�9z*�9�)�9�)�9(*�9,�9�+�9�+�9,�9;*�9�*�9-,�9�'�9�)�9-�9D*�98*�9x   x   �)�9�)�9�,�9+�9(+�9�'�9�*�9�/�9�-�9a+�9B0�9]+�9\-�9(/�9*�9)�9e,�9p*�9f-�9�(�9"*�9}.�9+�9M(�9 *�9�'�9�'�9e(�9�+�9�-�9x   x   �(�9_,�9!*�9^*�93+�9,�9�,�9�)�9Q&�9�)�9`+�9/&�9s*�9�-�92+�9*�9%)�9�*�9,�9)�9,�9�-�9q,�9�)�9,�9 -�9�+�9,+�9�-�90-�9x   x   �*�9f,�9-�9�'�9s*�9�,�9n(�9*�9�.�9�/�9[-�9r*�9�&�98-�9K+�9})�9.�9�*�9+�9,-�9Z*�9g*�9,�9x,�9�(�9+�9�+�9�+�9�)�9�,�9x   x   �'�9-(�9�-�9�'�9�,�9�,�9�,�9F.�9�+�9,�9+/�9�-�95-�9,�9&�9�+�9�(�9D)�9�,�9)�9�*�9�(�9�(�9�*�9�+�9-)�9�(�91*�9Y)�93.�9x   x   �(�9�(�9�*�9�%�9�+�9+�9�,�9;*�9�&�9|*�9!*�98+�9L+�9~&�9�,�9])�9K'�9F.�9E+�9�,�9--�9�,�9�+�9Z.�9�+�9�,�9h,�9.�9p)�9�.�9x   x   �&�9�*�9�-�9�(�9S*�9�'�9J(�9r,�94+�9�)�9)�9*�9z)�9�+�9`)�9)'�9:+�9l&�9�(�9�*�9�+�9�,�9�,�9�+�9Y,�9�,�99*�9�(�9&'�9g*�9x   x   �&�9'�9q-�9j)�9C-�9�*�92,�9�.�9�+�9�)�9h,�9")�9.�9�(�9N'�98+�9^,�9�+�9})�9�+�9=,�9R,�9
)�9.�9L+�9,�9 )�93,�9,�9u+�9x   x   �*�9�*�9�+�9)�9R)�9�+�9(�9w)�9�+�9**�9m*�9�*�9�*�9F)�9J.�9k&�9�+�9#,�9-�9c+�9�,�9�/�9x-�9�,�9�+�9�-�9�+�9�*�9Z'�9s.�9x   x   �*�9�+�9i-�9�-�9B-�9W,�9�'�95+�9).�9,�9d-�9,�9+�9�,�9@+�9�(�9�)�9-�9�,�9+�9�'�9g)�9&)�9�+�9�+�9-�9�*�9�(�9�)�9�+�9x   x   p)�9)�9�*�9-�9m,�9�*�9�*�9�,�9V-�9�+�9�(�9)�9*-�9)�9�,�9�*�9�+�9d+�9+�9\/�9'+�9�+�9\-�9M+�9C,�9�*�9*�97-�9�+�9�,�9x   x   �)�9�,�9m)�9,+�9�,�9r(�9�,�9�)�9�)�9�+�9#*�9,�9W*�9�*�9.-�9�+�9;,�9�,�9�'�9'+�9F+�9^+�9�)�9	,�9+,�9�,�9�-�9(�9)�9�,�9x   x   w+�9�-�9U*�9�-�9�+�9�*�9}.�9�*�9T-�9,�9�.�9�-�9f*�9�(�9�,�9�,�9Q,�9�/�9g)�9�+�9]+�9�(�9.�9 -�9�,�9+�9�*�9m,�9.�9&.�9x   x   �+�9,�9�*�9�)�9L,�9K)�9*�9�+�9U,�9:*�9+�9u,�9~,�9�(�9�+�9~,�9)�9{-�9$)�9\-�9�)�9.�9^*�9Y+�9z-�9l(�9+*�9�+�9�*�9�+�9x   x   t+�9J,�9)�9�+�9�,�9)�9�,�9�*�9�+�9�*�9M(�9�)�9u,�9�*�9X.�9�+�9.�9�,�9�+�9L+�9,�9"-�9Y+�94.�9�*�9�-�9�*�9�)�9Z)�9.+�9x   x   +�9�(�9$+�9�,�9K*�9�(�9H+�9�(�9�*�9.,�9*�9,�9�(�9�+�9�+�9Z,�9M+�9�+�9�+�9D,�9-,�9�,�9y-�9�*�9"(�9,�9�'�9�,�9�+�9�(�9x   x   �)�9�'�9�(�9�(�9F)�9)�9&,�9�'�9�,�9�'�9�'�9$-�9+�9/)�9�,�9�,�9,�9�-�9-�9�*�9�,�9+�9m(�9�-�9,�97)�9�(�9�+�9�'�9,�9x   x   �,�9s+�9w*�9�*�9,�9i-�93-�9�)�9-�9�)�9�'�9�+�9�+�9�(�9i,�9<*�9$)�9�+�9�*�9*�9�-�9�*�9&*�9�*�9�'�9�(�9�,�9]*�9�-�9�,�9x   x   -�9t,�9=-�91-�9�*�9*(�9e-�9�)�9|+�9-�9f(�90+�9�+�90*�9.�9�(�94,�9�*�9�(�97-�9(�9p,�9�+�9�)�9�,�9�+�9]*�9g,�9(�9�*�9x   x   �*�9�.�9*�9�/�9B,�9Z'�9�-�9�(�9�*�9B*�9�+�9�-�9�)�9Y)�9k)�9&'�9	,�9['�9�)�9�+�9)�9.�9�*�9Y)�9�+�9�'�9�-�9(�9�,�9/�9x   x   ,�9�,�9Z%�9�.�9/,�9 -�9R+�9%)�9�+�96*�9�-�9.-�9�,�91.�9�.�9g*�9v+�9r.�9�+�9�,�9�,�9.�9�+�9-+�9�(�9,�9�,�9�*�9/�9L%�9x   x   �;�9Z?�9U=�9_;�9*=�9�=�9@�9�;�9Y=�9+=�9m>�92>�9+=�9�=�9~?�9�>�9J>�9=@�9E=�9f>�9J>�9�;�9�=�9�<�9�?�9�<�9>�9�;�98=�9W?�9x   x   W?�9�;�9�;�9^A�9@�9cA�95=�9�=�9�=�9c?�9JD�9�<�9�?�9E�9Y@�9�A�9�C�92>�9�<�9�D�9F@�9�=�9#=�9<�9fB�9�@�99@�9;�9<�9d?�9x   x   T=�9�;�9hA�9�?�9;B�9j?�97>�9QB�9Q<�9<�9�A�9�:�95>�9�>�9�;�9+?�94?�9|<�9�@�9�:�9�<�9CB�9'?�9�?�9�@�9�?�9C�9�;�9�<�9r?�9x   x   ^;�9aA�9�?�9�8�9'<�9�?�9n<�9?�9 <�9E<�9�@�9�>�9D>�9�B�9�@�9�>�9�=�9I?�9>>�9e<�9�>�9<�9H?�9"<�9�9�9%?�9�?�9�;�9H=�9R<�9x   x   *=�9	@�97B�9%<�9�@�9�>�9�9�9y>�9�>�9�<�93=�9#A�9�>�9�?�9C@�9�@�9�>�9�<�9�=�9>�9�:�9?�9A�9
<�9XA�9-A�9i>�9�>�9x?�9�?�9x   x   �=�9iA�9g?�9�?�9�>�9	@�9�A�9�<�9�>�9�@�9�>�9>=�9�;�9~;�9<<�9X?�9�?�9V>�9k>�9iA�9>?�9�>�9P?�9�?�9B�9M<�9b=�9�=�9=�9�=�9x   x   @�96=�96>�9k<�9�9�9�A�9�A�9�?�9�;�9�?�9n?�9o>�9�C�9�>�9h@�9�>�9�=�9?�9�@�9dB�9�9�9�<�9�>�9�<�9 @�9.?�9�>�9�?�9�>�9�=�9x   x   �;�9�=�9UB�9?�9z>�9�<�9�?�9]?�9�<�9�B�9<�9k=�9�=�9f;�9�B�9�<�9�=�9�?�9G=�9�>�9w>�9�A�9y=�9�;�9B�9b?�9�=�9�=�9�@�9B�9x   x   Z=�9�=�9R<�9!<�9�>�9�>�9�;�9�<�9C�9;�9}<�9#A�9�<�9�:�9�C�9#<�9g=�9�>�9�=�9g<�9=�9�=�9	>�9m@�9@?�9�=�9�?�9!<�9D?�9�@�9x   x   *=�9a?�9<�9G<�9�<�9�@�9�?�9�B�9;�9U;�9�?�9<?�9�;�9�:�9�B�9�?�9$>�9�=�9�<�9�;�9?�9V<�9]>�9�=�9?�9
@�9B�9�?�9�<�9�>�9x   x   n>�9MD�9�A�9�@�95=�9�>�9s?�9<�9}<�9�?�9�8�9�?�9�<�9�;�9�>�9G@�9�>�9~?�9kA�9D�9p?�9�=�9�<�9+>�9OC�9�=�9]A�9�>�9\=�9�<�9x   x   3>�9�<�9�:�9�>�9"A�9@=�9r>�9k=�9%A�97?�9�?�9�@�9>�9~?�9?<�9@�9�=�9�;�9V=�9�=�9D;�9�>�9	=�9�>�9�<�9c=�9�?�9<�9!?�9�<�9x   x   '=�9�?�9/>�9A>�9�>�9�;�9�C�9�=�9�<�9�;�9�<�9>�9�A�90<�9�?�94?�9L?�9;>�9	=�9�?�9�?�9�@�9�=�9)@�9�?�9�?�9E=�9�A�9�>�9�>�9x   x   �=�9E�9�>�9�B�9�?�9�;�9�>�9a;�9�:�9�:�9�;�9}?�9/<�9q?�9�A�9�=�9@E�9?�9S?�9�<�9v>�9M@�9�<�9�A�9WA�9�<�9x@�9X>�9p=�9@�9x   x   �?�9\@�9<�9�@�9B@�9:<�9l@�9�B�9�C�9�B�9�>�9=<�9�?�9�A�9�=�9�@�9�>�9|>�9yA�9?<�9m>�9s@�9L:�9S<�9�:�9�@�9�=�9=�9@�9�>�9x   x   �>�9�A�9?�9�>�9�@�9R?�9�>�9�<�9%<�9�?�9E@�9@�98?�9�=�9�@�9?�9-@�9�<�9�@�9�>�9�;�9�=�9>>�9�=�9�<�9�<�9�>�9H@�9�=�9@�9x   x   P>�9�C�91?�9�=�9�>�9�?�9�=�9�=�9f=�9">�9�>�9�=�9O?�9>E�9�>�9,@�9RA�9?�9�@�9X?�9j<�9j?�9h;�9�@�9�;�9E?�9�@�9U?�9"@�9�@�9x   x   9@�91>�9�<�9J?�9�<�9R>�9?�9�?�9�>�9�=�9~?�9�;�9=>�9?�9{>�9�<�9?�9�<�9�;�9�>�9	@�9
=�9�;�9@�9�>�9�;�9�<�9%?�9|=�9�>�9x   x   E=�9�<�9�@�9D>�9�=�9j>�9�@�9G=�9�=�9�<�9kA�9S=�9
=�9Q?�9{A�9�@�9�@�9�;�9$=�9>�9�;�9T>�9N<�9s>�9%=�9b;�9�@�9A�9�?�9�>�9x   x   j>�9�D�9�:�9e<�9>�9iA�9aB�9�>�9f<�9�;�9D�9�=�9�?�9�<�9@<�9�>�9X?�9�>�9>�9m?�9�?�9t@�9>�9�=�9s?�9t?�9�=�9�<�9?�9�>�9x   x   H>�9F@�9�<�9�>�9�:�9A?�9�9�9v>�9=�9?�9o?�9C;�9�?�9u>�9j>�9�;�9j<�9@�9�;�9�?�9<�9@�9a=�9N?�9�;�9=�9�>�9><�9�>�9�;�9x   x   �;�9�=�9FB�9<�9	?�9�>�9�<�9�A�9�=�9V<�9�=�9�>�9�@�9L@�9n@�9�=�9l?�9=�9U>�9w@�9@�9e=�9'<�9�@�9�<�9�>�9�A�9�A�9_?�9�=�9x   x   �=�9#=�9'?�9E?�9A�9M?�9�>�9x=�9	>�9Y>�9�<�9=�9�=�9�<�9I:�9B>�9h;�9�;�9O<�9>�9a=�9)<�9*;�9�=�9&<�9<�9*<�9K<�9�;�93@�9x   x   �<�9<�9�?�9&<�9<�9�?�9�<�9�;�9m@�9�=�9)>�9�>�9*@�9�A�9W<�9�=�9�@�9@�9s>�9�=�9O?�9�@�9�=�9�;�9�@�9A�9�?�9�?�9V<�9?�9x   x   �?�9cB�9�@�9�9�9[A�9�A�9@�9B�9>?�9?�9NC�9�<�9�?�9YA�9�:�9�<�9�;�9�>�9)=�9x?�9�;�9�<�9)<�9�@�9 @�9]<�9�@�9�?�9�@�9�A�9x   x   �<�9�@�9�?�9$?�90A�9P<�93?�9d?�9�=�9
@�9�=�9c=�9�?�9�<�9�@�9�<�9C?�9�;�9b;�9s?�9=�9�>�9<�9A�9V<�9@�9�@�9<�9c?�9+?�9x   x   >�97@�9C�9�?�9h>�9a=�9�>�9�=�9�?�9	B�9\A�9�?�9G=�9v@�9~=�9�>�9�@�9�<�9�@�9�=�9�>�9�A�9*<�9�?�9�@�9�@�9�@�9>�9�>�9$=�9x   x   �;�9;�9�;�9�;�9�>�9�=�9�?�9�=�9<�9�?�9�>�9<�9�A�9W>�9=�9G@�9U?�9$?�9A�9�<�9><�9�A�9L<�9�?�9�?�9<�9>�9�>�9�=�9?�9x   x   5=�9<�9�<�9E=�9y?�9=�9�>�9�@�9E?�9�<�9Z=�9 ?�9�>�9w=�9 @�9�=�9"@�9|=�9 @�9?�9�>�9_?�9�;�9X<�9�@�9b?�9?�9�=�9.?�9�<�9x   x   W?�9g?�9p?�9S<�9�?�9�=�9�=�9B�9�@�9�>�9�<�9�<�9�>�9@�9�>�9@�9�@�9�>�9>�9�>�9�;�9�=�93@�9?�9�A�9'?�9%=�9?�9�<�9?�9x   x   	N�9HR�9sY�9�T�9T�9�U�9�T�9�S�9�U�9�S�9�S�9KU�9V�9hR�9�S�9�T�9�R�9�R�9�V�9?U�9�S�9�R�9*V�9�U�9�S�9sT�9�T�9?U�9�Y�9FR�9x   x   IR�9�S�9�U�9�Q�9�P�9�O�9�T�9�U�9uQ�9�S�9~O�9-S�9/U�9xO�9�R�9�S�9�O�9]T�9�R�9$P�9RT�9�Q�9�T�9WS�9fQ�9�Q�9�P�9DU�9�S�9R�9x   x   sY�9�U�9P�9�R�9T�9�R�9�S�9�P�9�V�9�S�9�O�9�T�9�P�9.O�9DR�9�N�9LQ�9�U�9�O�9S�9�V�9'Q�9U�9�R�9AR�9�R�9�Q�9�U�9MY�9X�9x   x   �T�9�Q�9�R�9�V�9U�9AU�9�R�9�V�9�V�9�S�92V�9�V�9�S�9vU�9&U�9�S�9V�9�U�9�T�9W�9'V�9�Q�9�T�9}U�9kX�94R�9�P�9�T�9�Q�9-Q�9x   x   T�9�P�9T�9U�9�O�9�S�9KU�9NS�9�S�9|T�9ZP�9�S�9R�9P�9�R�9CS�9�P�9�T�98S�91S�9�V�9sS�9�O�9�T�9
S�9{Q�9PU�9/T�9cS�9�T�9x   x   �U�9�O�9�R�9BU�9�S�9|V�9kP�9Q�9�T�9�U�9�S�9*U�9T�9�S�9�T�9�T�9U�9�T�9�Q�9~O�9V�9T�9�T�9�R�9�P�9PT�9$T�9YV�9�U�9�T�9x   x   �T�9�T�9�S�9�R�9IU�9nP�9�R�9�T�9S�9�S�9R�9�R�9�T�9$S�9�Q�9�S�9T�9/T�9$S�9�P�9 U�9mR�9�T�9T�92T�9Q�9�Q�9�R�9�Q�9&P�9x   x   �S�9�U�9�P�9�V�9LS�9Q�9}T�9�U�9JR�9�P�9�R�9�S�9�S�9�R�9�P�9MR�9U�9�S�9!Q�9�S�9�V�9mP�9U�9VT�9Q�9'U�9]T�9�T�9�U�9�P�9x   x   �U�9tQ�9�V�9�V�9�S�9�T�9S�9LR�9?T�9fV�9V�9�U�9�U�9�V�9BT�9�Q�9�T�9*U�98S�9mV�9�V�9�Q�9VV�9YQ�9DR�9LS�9+S�9R�9�R�9!R�9x   x   �S�9�S�9�S�9�S�9|T�9�U�9�S�9�P�9fV�9�T�9mS�9�S�9uT�9�U�9�Q�9_S�9tT�9$U�9�T�9�S�9�S�9S�9�T�9U�9�P�9�P�9R�9(Q�9�S�9<U�9x   x   �S�9O�9�O�90V�9ZP�9�S�9R�9�R�9�U�9lS�9�Q�9S�9�V�9JR�9�Q�9	U�9Q�9U�9�O�9�O�9�T�9�T�9}V�9BV�9�R�9U�9�Q�9=W�9�V�9T�9x   x   HU�9)S�9�T�9�V�9�S�9+U�9�R�9�S�9�U�9�S�9�S�9�T�9�S�9HS�9�T�9�R�9�V�9xU�9S�9�T�9�S�9�P�9�T�9S�9�S�97T�9�R�99T�9�P�9�T�9x   x   V�9/U�9�P�9�S�9R�9T�9�T�9�S�9�U�9uT�9�V�9�S�9^T�9�S�9�R�9T�9�P�9�T�9�V�9�T�98T�9�P�9�S�9aR�9P�9�R�9�S�9^Q�9�S�9�S�9x   x   jR�9tO�9-O�9uU�9P�9�S�9#S�9�R�9�V�9�U�9KR�9LS�9�S�9P�9�T�9�N�9�O�9�R�9�O�9(T�9�U�9�R�9CV�9�R�9�Q�9V�9�R�9KU�9�T�9�P�9x   x   �S�9�R�9FR�9'U�9�R�9�T�9�Q�9�P�9>T�9�Q�9�Q�9�T�9�R�9�T�9�R�9�R�9lS�9�Q�9~T�9�S�9�Q�9yT�9#U�9&S�9�U�9pT�9�Q�95T�9sS�9eQ�9x   x   �T�9�S�9�N�9�S�9BS�9�T�9�S�9MR�9�Q�9aS�9U�9�R�9T�9�N�9�R�9U�9�R�9�S�9
T�9HS�9*U�9�T�9�V�9�V�9?T�9�U�9S�9T�9 U�9sR�9x   x   �R�9�O�9MQ�9�U�9�P�9U�9	T�9U�9�T�9tT�9
Q�9�V�9�P�9�O�9nS�9�R�9KR�9R�9IR�9�T�9�R�9^R�9YU�9�R�9�R�9�T�9tR�9�Q�9�Q�9>S�9x   x   �R�9^T�9�U�9�U�9�T�9�T�9-T�9�S�9,U�9!U�9!U�9vU�9�T�9�R�9�Q�9�S�9R�9[U�9lU�9~S�9�R�9U�9�T�9�R�9jS�9�U�9�U�9ER�9�S�9 R�9x   x   �V�9�R�9�O�9�T�97S�9�Q�9'S�9#Q�9:S�9�T�9�O�9S�9�V�9�O�9~T�9T�9HR�9oU�9eU�9nT�97U�9�X�9wU�9�T�9uU�9�T�9;R�9�T�9~S�9�O�9x   x   >U�9%P�9S�9W�9.S�9�O�9�P�9�S�9jV�9�S�9�O�9�T�9�T�9#T�9�S�9FS�9�T�9�S�9nT�9�R�9S�9/S�9/R�94T�9T�9�U�9%R�9OT�9+U�9�S�9x   x   �S�9TT�9�V�9(V�9�V�9�U�9�T�9�V�9�V�9�S�9�T�9�S�99T�9�U�9�Q�9+U�9�R�9�R�98U�9S�9�O�9.S�9�U�9:R�9�Q�9/V�9*R�9�T�9#T�9T�9x   x   �R�9�Q�9'Q�9�Q�9xS�9!T�9oR�9lP�9�Q�9S�9�T�9�P�9�P�9�R�9{T�9�T�9\R�9U�9�X�9*S�9+S�9/X�9�T�9�S�9�S�9�S�92S�9OQ�9Q�9�T�9x   x   .V�9�T�9�T�9�T�9�O�9�T�9�T�9U�9SV�9�T�9|V�9�T�9�S�9EV�9U�9�V�9[U�9�T�9yU�9.R�9�U�9�T�9T�9�V�9<V�9V�9yS�9]T�9�U�9�U�9x   x   �U�9WS�9�R�9}U�9�T�9�R�9T�9WT�9\Q�9 U�9FV�9S�9`R�9�R�9"S�9�V�9�R�9�R�9�T�94T�99R�9�S�9�V�9�R�9%R�9�R�9�S�9|W�9AT�9oP�9x   x   �S�9fQ�9@R�9gX�9S�9�P�90T�9Q�9ER�9�P�9�R�9�S�9P�9�Q�9�U�9?T�9�R�9iS�9rU�9T�9�Q�9 T�9:V�9%R�9�P�9�S�9�P�9_Q�9�S�9�P�9x   x   mT�9�Q�9�R�92R�9~Q�9OT�9 Q�9(U�9KS�9�P�9U�94T�9�R�9V�9oT�9�U�9�T�9�U�9�T�9�U�91V�9�S�9V�9�R�9�S�9�V�9Q�9�Q�9KU�9*Q�9x   x   �T�9�P�9�Q�9�P�9OU�9 T�9�Q�9]T�9*S�9R�9�Q�9�R�9�S�9�R�9�Q�9S�9rR�9�U�9<R�9'R�9*R�93S�9{S�9�S�9�P�9Q�9T�9�T�9�Q�95T�9x   x   >U�9@U�9�U�9�T�92T�9YV�9�R�9�T�9R�9*Q�9<W�96T�9cQ�9LU�92T�9T�9�Q�9FR�9�T�9MT�9�T�9QQ�9\T�9wW�9_Q�9�Q�9�T�9qR�9:V�9�T�9x   x   �Y�9�S�9LY�9�Q�9eS�9�U�9�Q�9�U�9�R�9�S�9�V�9�P�9�S�9�T�9sS�9�T�9�Q�9�S�9~S�9+U�9 T�9Q�9�U�9=T�9�S�9KU�9�Q�99V�9%S�9nQ�9x   x   FR�9R�9X�9*Q�9�T�9�T�9#P�9�P�9 R�9>U�9T�9�T�9�S�9P�9hQ�9sR�9=S�9 R�9�O�9�S�9T�9�T�9�U�9mP�9�P�9(Q�94T�9�T�9nQ�9�W�9x   x   �x�9�i�9�e�9Ui�9=i�9�k�9k�9{i�9wi�9Rj�9Ui�9Gh�9�g�9<l�9*k�9 g�9 j�9�j�9�h�9�g�9�i�9cj�9-i�9�j�9sj�9�j�9�i�9xi�9�e�9�i�9x   x   �i�9�f�9ti�9k�9*k�9�h�9Kj�9j�9vj�9[j�9i�9�l�9Th�9�i�9bj�9�j�9gk�9�h�94l�9�h�9$j�9?k�9�h�9�i�9/j�9#k�9�j�9�i�9�f�9�i�9x   x   �e�9ri�9Fj�9�j�9�h�9�h�9�i�9h�9wh�9�l�9	k�9j�9m�9�o�9`l�9�n�9�k�9�i�9Ml�9Am�9�g�9�h�9�j�9h�90h�9�j�9Wj�9Zi�9f�9�b�9x   x   Ui�9k�9�j�94h�9�i�9�j�9�j�9:f�9le�9k�9Mg�9�g�9�i�9mg�9�h�9�j�9�h�9
g�9�i�9qf�9�e�9tj�9�j�9�i�9�h�9�j�9k�9Hi�9k�9Nk�9x   x   @i�9,k�9�h�9�i�9�h�9i�9l�9�i�9i�9 i�9�i�9h�9-i�9j�9Ch�9�g�9i�9j�9�h�9j�9�l�9�h�9*i�9�i�9Uh�9?k�9Zi�9�g�9�j�9�g�9x   x   �k�9�h�9�h�9�j�9 i�9�f�9�i�9�n�9?h�9�g�9�h�9�j�9-n�9�m�9�k�9	i�9�g�9�h�9in�9�h�9Dg�9Wi�9Xj�9�h�9oi�9wk�9�i�9�g�9hg�9�i�9x   x   k�9Lj�9�i�9k�9l�9�i�9�k�9�f�9�h�9j�9�j�98i�9�c�9�i�9�i�9�j�9�g�9mf�9�l�9�i�9�k�9�j�9Hj�9�i�9�j�9�j�9k�9�h�9Uk�9�j�9x   x   |i�9j�9h�9<f�9�i�9�n�9�f�9j�9qm�9)h�9�n�9:j�9�i�9�n�9h�9�m�9k�9�e�9@n�9�i�9�f�9�g�9�i�9j�9�i�9�i�9.i�9i�9�i�9Ni�9x   x   si�9yj�9wh�9je�9i�9Bh�9�h�9wm�9�e�9i�9�g�9�c�9�g�9�i�9%e�9 m�9�h�9�h�9�i�9e�94h�9�j�9�i�9Zi�9�k�9k�9fj�9�j�9(l�9
j�9x   x   Rj�9]j�9�l�9k�9i�9�g�9j�9*h�9i�9i�9eh�9Ai�9�g�9�h�9wi�9gi�96h�9�h�9k�9�l�9<j�9j�9�f�9�i�9�l�9�k�9�k�9�l�9�h�9�f�9x   x   Vi�9i�9	k�9Og�9�i�9�h�9�j�9�n�9�g�9nh�9�q�9�h�9Ni�9�m�9uj�9Oi�9Si�9�f�9Xk�9�i�9+i�9(j�9&f�9"f�9g�9�i�9�f�9�f�9�f�9j�9x   x   Gh�9�l�9j�9�g�9h�9�j�99i�9?j�9�c�9Gi�9�h�9@c�9|i�9�i�9 k�9,g�9,i�9�j�9�k�9�g�9�k�9�k�9�k�9zh�9rl�9�l�9�g�9 k�9�k�9ck�9x   x   �g�9Vh�9m�9�i�9/i�9-n�9�c�9�i�9�g�9�g�9Gi�9wi�9�d�9fm�9�i�9�i�9Vk�9�h�9�h�9�g�9�h�9�i�9ek�9�i�97l�9�i�9�k�9�i�9�i�9[g�9x   x   <l�9�i�9�o�9jg�9 j�9�m�9�i�9�n�9�i�9�h�9�m�9�i�9fm�9Vj�9�g�9�p�9=j�9sk�9�k�9�i�9�j�9�h�9i�9gj�9�i�9�h�9_h�9�i�9�i�9�l�9x   x   *k�9hj�9[l�9�h�9Ch�9�k�9�i�9h�9$e�9yi�9vj�9 k�9�i�9�g�9k�9wj�9�j�9ym�9*h�9�i�9�j�9ef�9�i�9�i�9lj�9f�9vk�9�i�9�g�9�l�9x   x   g�9�j�9�n�9�j�9�g�9i�9�j�9�m�9 m�9ei�9Mi�9+g�9�i�9�p�9tj�9�f�93i�9�j�90h�9�j�9k�9xh�9vf�9#f�9sh�9�j�9j�9�h�9�k�9�h�9x   x   �i�9ck�9�k�9�h�9i�9�g�9�g�9k�9�h�95h�9Si�9,i�9Xk�9:j�9�j�93i�9|j�9k�9�f�9"h�9�l�9i�9�i�9�h�9m�9�g�9�f�9,j�9k�9�i�9x   x   �j�9�h�9�i�9g�9j�9�h�9kf�9�e�9�h�9�h�9�f�9�j�9�h�9rk�9ym�9�j�9k�9Gl�9Bi�9ih�9�j�9�h�9i�9j�9rh�9�i�9�l�9�j�9Cj�9�m�9x   x   �h�95l�9Ml�9�i�9�h�9dn�9�l�9:n�9�i�9k�9Vk�9�k�9�h�9�k�9+h�90h�9�f�9Ai�9Ah�9ci�9�h�9bc�9�h�9ii�9�g�9xh�9/g�9�h�9�g�9�l�9x   x   �g�9�h�9Am�9tf�9j�9�h�9�i�9�i�9e�9�l�9�i�9�g�9�g�9�i�9�i�9�j�9 h�9eh�9^i�9�i�9-i�9�h�9aj�9�i�9i�9dh�9�i�9wj�9�h�9�g�9x   x   �i�9!j�9�g�9�e�9�l�9Bg�9�k�9�f�91h�96j�9+i�9�k�9�h�9�j�9�j�9k�9�l�9�j�9�h�91i�9�q�94i�9=h�9:j�9�k�9�k�9�j�9�j�9bi�9�k�9x   x   ej�9@k�9�h�9sj�9�h�9Yi�9�j�9�g�9�j�9j�9*j�9�k�9�i�9|h�9ff�9{h�9�h�9�h�9bc�9�h�96i�9yc�9Ci�9�i�9#h�9kf�9�g�9�i�9uk�9�i�9x   x   ,i�9i�9�j�9�j�9)i�9]j�9Ij�9�i�9�i�9�f�9(f�9�k�9ak�9i�9�i�9xf�9�i�9i�9�h�9bj�9;h�9Ci�9Nh�9�f�9�i�9vi�9�k�9Ok�9g�9�f�9x   x   �j�9�i�9h�9�i�9�i�9�h�9�i�9j�9Xi�9�i�9 f�9yh�9�i�9fj�9�i�9$f�9�h�9j�9ii�9�i�99j�9�i�9�f�9�i�9.j�9i�9|h�9�e�9Hi�9�i�9x   x   uj�90j�90h�9�h�9Th�9ri�9�j�9�i�9�k�9�l�9g�9sl�98l�9�i�9rj�9sh�9m�9rh�9�g�9#i�9�k�9 h�9�i�9/j�9�l�9�l�9�g�9�l�9�k�9�h�9x   x   �j�9#k�9�j�9�j�9;k�9xk�9�j�9�i�9k�9�k�9�i�9�l�9�i�9�h�9f�9�j�9�g�9�i�9xh�9fh�9�k�9kf�9wi�9i�9�l�9�h�9�k�9k�9j�9^k�9x   x   �i�9�j�9Wj�9k�9\i�9�i�9k�90i�9gj�9�k�9�f�9�g�9�k�9Zh�9sk�9~j�9�f�9�l�9.g�9�i�9�j�9�g�9�k�9|h�9�g�9�k�9Xj�9i�9�j�9j�9x   x   yi�9�i�9\i�9Ii�9�g�9�g�9�h�9i�9�j�9�l�9�f�9 k�9�i�9�i�9�i�9�h�9/j�9�j�9�h�9wj�9�j�9�i�9Qk�9�e�9�l�9k�9 i�9�i�9Kg�9Cg�9x   x   �e�9�f�9f�9k�9|j�9hg�9Sk�9�i�9'l�9�h�9�f�9�k�9�i�9�i�9�g�9�k�9k�9Bj�9�g�9�h�9bi�9vk�9g�9Ii�9�k�9j�9�j�9Ng�9!k�9k�9x   x   �i�9�i�9�b�9Pk�9�g�9�i�9�j�9Pi�9j�9�f�9j�9ek�9_g�9�l�9�l�9�h�9�i�9�m�9�l�9�g�9�k�9�i�9�f�9�i�9�h�9ak�9j�9Hg�9k�9�b�9x   x   �u�9���9���9Ҁ�9��9�|�9��9��9��9o��98��9��9�~�9���9W��9x��9ۀ�9K~�9/�9Q��9^��9h��9�~�9j��9�~�9�|�9ހ�9ƀ�9c��9��9x   x   ���9���9e��9���9��9���9���9H�9B��9��9���9��9 �9*��9��9L�9w��9��9��9ց�9y~�9���9�~�9n��9���9��9���9��9���9��9x   x   ���9h��97��9��9'��9��9���9Ć�9Q��9��9���9%��9̀�9��9&}�98~�9j�9�~�9���9���9���9���9#��9���9��9N��9��9��9ӂ�9*��9x   x   Ӏ�9���9߀�9�~�9��9m�9���9D��91��9���9a��9��9��9���9���9e��9ȁ�9w��9��9-��9���9���9A��9��9�}�9%��9n��9��9���9���9x   x   ��9��9#��9��9���9���9��9���9���9V��9w��9Z��9'��9���9���9��9Z��9v��9Y��9��9��9��9z��9��9ۃ�9	��9��9��9=��9t��9x   x   �|�9���9}��9q�9���9���9r��9��9���9<��9���9�}�9�~�9�~�9[�9���9��9o��9_�9=��9��9ہ�9��9E��9T��9~�9{��9+��9���9���9x   x   ��9���9���9���9��9q��9�9k��9���9=��9���9��9��9��9 ��9ł�9��9���9��9*��9��98��9р�9e��9A�9Ѐ�9���9��9
��9���9x   x   ��9L�9���9C��9���9��9l��9�~�9�9���9�}�9��9���9f~�9ł�9	�9(��9��9��9s��9���9���9d�9���9���9-�9���9���9V~�9Ƀ�9x   x   ��9D��9Q��91��9���9���9���9�9��9���9�~�9��9�~�9ā�9'��9�~�9���9���9��9���9s��9O��9�~�9���9�~�9i}�9}��9�~�9y~�9(��9x   x   m��9��9��9���9V��98��9?��9���9���9���9��9��9o��9m��9��9���9���9���9���9o�9]�99��9���9U��9Ɓ�9���9���9���9W��9?��9x   x   6��9���9���9e��9x��9���9���9�}�9�~�9��9�x�9��9'��9~}�9ـ�9���9���9[��9���9G��9l��9��9]��9ł�9 ��9k~�9p��9Ղ�9���9L��9x   x   	��9��9&��9 ��9]��9�}�9��9��9݆�9��9��9���97��9��9�~�9׃�9ˁ�9��9Y��9��9���9 ��9p��9؃�9d~�9�~�9F��9{��9ǁ�9��9x   x   �~�9�~�9ɀ�9��9!��9�~�9	��9���9�~�9v��9/��9<��9'��9�}�9��9x�9,�9(��9�~�9��9Z��94��9��9U��9���9��9���9���9-��98��9x   x   ���9(��9��9���9���9�~�9��9g~�9Ɓ�9l��9~}�9��9�}�9���9k��9q��9���9��9���9ǂ�9��9؄�9L��9<��98��9k��9���9��9���9|��9x   x   W��9��9'}�9���9���9Y�9��9Â�9)��9��9׀�9�~�9��9j��9�{�9��9���9�}�9��9��9ȁ�9���9���9���9
��9*��9���9J�9%��9}�9x   x   s��9J�9:~�9f��9��9���9ǂ�9�9�~�9��9���9׃�9z�9o��9��9���9F��9���9F��9҂�9�}�9#��9���9G��9���9�}�9ł�9���9���9́�9x   x   ݀�9v��9g�9΁�9X��9
��9��9 ��9���9���9���9́�9-�9���9À�9G��9b��9���9J��9��9���9��96��9���9��9���9z��9��9���9P��9x   x   N~�9��9�~�9x��9v��9p��9���9��9���9���9X��9��9'��9��9�}�9���9���9�~�9���9t��9���9΁�9���9.��9҂�9ށ�9@�9���9��9~�9x   x   +�9��9���9��9Z��9_�9��9��9��9���9���9Y��9�~�9���9��9E��9F��9���9͂�9��9j��9_��9'��9Հ�9���9 ��9g��9���9��9���9x   x   Q��9Ձ�9���9+��9��9=��9+��9t��9���9t�9G��9��9��9ǂ�9��9Ԃ�9��9x��9	��9ρ�9���9��9�9���9 ��91��9c��9+��9΀�9v��9x   x   [��9y~�9���9���9��9��9��9���9p��9_�9m��9���9\��9��9ȁ�9�}�9���9���9i��9���9�9���9���9u��9��97~�9~��9��93��9:��9x   x   g��9���9���9���9��9ځ�97��9���9O��99��9��9���95��9ۄ�9���9 ��9��9΁�9^��9
��9���9o��9���9P��9T��9#��9���9l��9���9�~�9x   x   �~�9�~�9%��9E��9|��9��9π�9d�9�~�9���9_��9s��9��9J��9݂�9���98��9���9&��9���9���9���9��9ׂ�9���9>��9��9���9��9���9x   x   i��9i��9���9��9��9E��9b��9���9��9V��9Ƃ�9ڃ�9Y��9;��9���9F��9���9/��9׀�9���9s��9Q��9ق�9J��9T��9�~�9h��9��9ނ�9��9x   x   �~�9���9��9�}�9܃�9T��9A�9���9�~�9ˁ�9���9a~�9���95��9��9���9��9҂�9���9��9��9Q��9���9R��9@��9�9��9a��9~�9��9x   x   �|�9��9N��9)��9	��9~�9Ѐ�9*�9j}�9���9l~�9�~�9��9m��9)��9�}�9���9߁�9!��9-��97~�9(��9@��9�~�9�9�{�9���9?~�9��9
��9x   x   ܀�9���9��9o��9��9}��9���9���9}��9���9m��9G��9���9���9���9ł�9v��9A�9j��9a��9��9���9��9g��9��9���9��9��9&��9��9x   x   ƀ�9��9��9���9��9,��9���9���9�~�9���9ւ�9~��9��9��9K�9���9��9���9���9.��9��9j��9���9��9a��9?~�9��9ڄ�9��9��9x   x   `��9���9ς�9���9?��9���9��9T~�9x~�9Y��9���9ǁ�9+��9���9"��9���9���9��9��9ʀ�93��9���9
��9܂�9~�9��9&��9��9,��9!��9x   x   ��9��9(��9��9s��9���9���9ȃ�9(��9<��9L��9��94��9{��9}�9́�9Q��9~�9���9q��98��9�~�9���9��9��9��9��9��9!��9���9x   x   ��9��9��9���9̝�9���9���9��9���9��9b��9��9��9���9���9��9i��9���98��9��9Y��9��9ƚ�9���9g��9���9���9p��9���9ٛ�9x   x   ��9��9��9Ę�9&��9��9��9��9��9��9���9��9i��9;��9)��9��9e��9��9~��9���9���9ژ�9p��9���9&��9���9Ǚ�9Ԛ�90��9̛�9x   x   ��9��9:��9_��9���9��9S��9���9���9N��9��9Ǟ�9A��9���9;��9$��9���9v��9E��9��9&��9���9b��9B��9���9��9��9��9S��9A��9x   x   ���9Ƙ�9a��9#��9��9��9ә�9u��9���9���9��9o��9���9Û�9d��9x��9���9���9���9��9(��9Y��9���9f��9u��9ə�9��9m��9���9��9x   x   ǝ�9'��9���9��9%��9���9���9���9r��9���9��9��9���9��9���9��9O��9���9���9C��9ݘ�9\��9���9-��9��9x��9@��9���9��9ʚ�9x   x   ���9��9��9���9���9m��9��9L��9���9���9���9)��9��9���9h��9ǘ�9���9Κ�9X��9F��9��9.��9��9h��9���9���9N��9���9���9��9x   x   ���9��9R��9ҙ�9���9��9���9���9Μ�9��9D��9���9I��9p��9ɛ�9ʚ�9���9B��9���9���9��9���9���9Κ�9���9���9���9��9���9��9x   x   ��9��9���9t��9���9K��9ě�9���9\��9g��9���9k��9���9���9%��9��9���9���93��9ܚ�9&��9j��9���9���9���9	��9/��9ԛ�9"��9��9x   x   ���9��9���9���9o��9���9ќ�9T��9���9��9���9��9n��9���9���9���9���9˚�9x��9���9���9���9���9ݖ�9��9r��9���9��9,��9���9x   x   ��9��9Q��9���9���9�9���9i��9��9u��9���9ϛ�9���9��9���9���9��9r��9D��9���9���9A��9,��9��9V��9x��9���9F��9��9͙�9x   x   f��9���9��9��9}��9���9B��9���9���9���9f��9���9��9���9��9��9���9-��9G��9 ��9���9��9k��9;��9��9R��9V��9���9ޛ�9m��9x   x   ��9��9ʞ�9m��9��9.��9���9f��9��9Λ�9���9��96��9���9כ�9Q��9_��9��9ܗ�9��95��9���9̗�9���9͙�9���9ٙ�9Ø�9���9m��9x   x   ��9k��9G��9���9���9��9F��9���9k��9���9��94��9���9���9��9��9���9p��9_��9_��9(��9��9!��9D��9���9��9���9(��9���9���9x   x   ���9<��9���9���9��9���9r��9���9���9��9���9���9���9>��9���9\��9��9J��9��9}��9r��9���9~��9͙�9&��9ٙ�9b��9)��9T��9+��9x   x   ���9)��9:��9b��9���9l��9ț�9&��9���9���9��9؛�9��9���9C��9͛�9���9���9���9��9%��9���9��9��9���92��9���9���9ĝ�9ܙ�9x   x   ��9��9&��9t��9��9ǘ�9Κ�9��9���9���9��9N��9��9_��9˛�9m��9���9+��9��9g��9��9���9ę�9��9��9ݚ�9��9���9K��91��9x   x   h��9g��9���9���9M��9Ŗ�9���9���9���9��9���9]��9��9��9���9���9x��9i��9ә�9m��9��9���9V��9��9ߚ�9��9���9��9G��9���9x   x   ���9��9t��9���9���9ǚ�9@��9���9Ț�9q��90��9��9l��9K��9���9-��9g��9=��9���9ؚ�9���9��9!��9���9���9ט�9t��9���9���9.��9x   x   6��9���9F��9���9���9Z��9���96��9{��9E��9I��9��9b��9��9���9��9ԙ�9���9���9��9q��9��9ә�9h��9��9p��99��9M��9ۜ�9���9x   x   ���9���9��9��9@��9B��9���9ۚ�9���9���9��9��9]��9{��9��9g��9l��9֚�9��9Ζ�9���9[��9��9Q��9��9��9���9���9Q��9ř�9x   x   [��9���9(��9)��9ܘ�9��9��9(��9���9���9���97��9(��9o��9$��9��9��9���9r��9���9u��9���9���9���9��9˚�9��9i��9R��9���9x   x   ��9֘�9���9X��9Z��9-��9���9l��9���9A��9~��9���9
��9���9���9���9���9��9��9W��9���9��9җ�9���9X��9V��9=��9X��9q��9j��9x   x   ɚ�9j��9c��9���9���9��9���9���9���9.��9j��9ɗ�9��9~��9��9�9S��9 ��9ؙ�9��9 ��9ӗ�9W��9*��9���9Z��9ښ�9���99��9Ϙ�9x   x   ���9���9F��9f��9,��9m��9Қ�9���9ݖ�9��98��9���9A��9ϙ�9��9��9��9���9j��9Q��9���9���9+��9���9H��9���9���9���9 ��9S��9x   x   f��9,��9���9q��9��9���9���9���9��9U��9 ��9Ι�9���9*��9���9���9ޚ�9���9��9��9#��9V��9���9I��9=��9���9��9$��9*��9:��9x   x   ��9���9��9ș�9z��9���9���9��9n��9t��9U��9���9��9י�94��9���9��9٘�9o��9��9Ϛ�9R��9W��9���9���9���9���9���9��9ɛ�9x   x   ���9ʙ�9|��9��9>��9J��9���93��9���9���9Z��9ڙ�9���9_��9���9��9���9u��9:��9���9���99��9���9���9��9���9՛�9���9ܔ�9ӛ�9x   x   n��9֚�9���9p��9���9���9��9כ�9��9D��9~��9���9'��9&��9���9���9��9��9L��9���9j��9V��9���9���9$��9���9�9���9ٚ�9`��9x   x   ���91��9T��9���9��9���9���9$��9*��9
��9ߛ�9���9���9S��9ǝ�9M��9D��9���9ۜ�9P��9W��9n��9:��9"��9,��9��9ܔ�9ۚ�9��9���9x   x   ڛ�9˛�9=��9	��9Ś�9ޚ�9��9��9���9Ι�9n��9o��9���9,��9��9/��9���92��9���9ƙ�9���9m��9Ϙ�9R��9>��9ƛ�9ϛ�9\��9��9���9x   x   y��9���9���9ٵ�9���9ʵ�9���9��9���9r��9���9E��9���9���9մ�9:��9w��9ͳ�9���9���9��9��9���9V��9��9*��9î�9���9���9���9x   x   ���9
��9=��9Z��9p��9b��9Ͳ�9���9r��9C��9���9���9���9(��9���9.��9��9A��9*��9u��9���9���9��9ճ�9��9Ҹ�9 ��9��9���9в�9x   x   ���9<��9b��9\��9���9���9���9g��9B��9���9��9���9���9���9���9J��9Y��9���9i��9y��9J��9���9G��9|��9ϲ�9���9��9���9<��9���9x   x   ۵�9Z��9X��9��9���9���9��9��9S��9���9X��9��9?��9���9��9��9Q��9x��9���9��9��9M��9:��9ε�9���9��9:��9��9/��9a��9x   x   ���9r��9���9���9ͱ�9 ��9
��9F��9]��9ܷ�9��9X��9���9g��9���9��9��9L��9��9��9��9���9��9δ�9���9���9%��9ĳ�9m��9ײ�9x   x   ȵ�9a��9���9���9!��9���9޳�9ն�9(��9V��9s��9��9 ��9 ��9)��96��9B��9$��9��9K��9��9��9���9��9���9���9԰�9z��9���9���9x   x   ���9в�9���9��9��9ݳ�9��9ñ�9.��9M��9α�9���9��9��9i��9���9W��9���9��9��9��9���9���9i��9���9:��9*��9η�9<��9U��9x   x   ��9���9k��9��9H��9׶�9ű�9���9���9d��9���9��9���9���9/��9r��9��9���9���9���9��9B��9#��9δ�9��9��9���9U��9���9<��9x   x   ���9p��9A��9P��9`��9"��9,��9���9��9o��9˹�9��9���9(��9Q��9>��9@��9���9��9:��9���9���9w��9 ��9ɷ�9u��9���9���9��9���9x   x   s��9A��9���9���9��9Q��9N��9g��9j��9���9���9K��9\��9г�9H��9���9��9���9��9��9f��9?��9���9���9'��9��9��9%��9շ�9��9x   x   ���9���9��9Y��9$��9p��9α�9���9ǹ�9���9��9���9���9V��9y��9���9���9���9&��9��9���9���9{��9���9���9���9V��9Ե�9F��9Y��9x   x   F��9���9���9��9Y��9��9���9��9��9O��9���9ʴ�9i��9��9ݲ�9v��9K��9ű�9	��9��9���93��9���9��9ѳ�97��9/��9���9X��9��9x   x   ���9���9��9<��9���9��9��9���9���9_��9���9c��9��9k��9A��9��9\��9l��9.��9v��9���9��9��9!��9���9v��9
��9j��92��9���9x   x   ���9#��9���9���9j��9��9��9���9)��9ӳ�9[��9��9k��9;��9/��9S��9���9p��9��9���9���9V��9A��9���9ȳ�9���9m��9���9���9��9x   x   Դ�9���9���9��9���9'��9j��93��9P��9K��9{��9ܲ�9C��9/��9���9��9���9���9'��9��9���9���9���9>��9��9Ѳ�9���9��9u��9��9x   x   ;��9/��9K��9��9��94��9���9l��99��9���9���9x��9��9S��9
��9���9��9׵�9-��9���9t��9A��9��9���9��9��9���9��9��9���9x   x   t��9��9\��9T��9��9?��9W��9$��9C��9��9���9N��9c��9���9���9��9���9q��9���9ѳ�9$��9Ͷ�9��9���9J��9W��9���9���9���9³�9x   x   γ�9>��9���9w��9N��9��9���9���9���9���9���9Ʊ�9j��9n��9���9յ�9r��9:��9���9���9���9?��9V��9��9,��9/��90��9��9���9]��9x   x   ���9,��9j��9���9��9��9��9���9��9��9%��9��9,��9��9%��9.��9���9���9���92��9���9��9��9���9
��9/��9���9g��9մ�9ڲ�9x   x   ���9q��9x��9��9��9M��9#��9���9=��9��9��9��9u��9���9��9���9г�9���93��9R��9���9���9���9 ��9���9[��9X��9���9��9���9x   x   ��9���9J��9��9��9��9��9��9���9f��9���9���9���9���9���9s��9'��9���9���9���9���9���9���9���9��9���9h��9���9���9(��9x   x   ��9���9���9K��9���9��9���9B��9���9?��9���94��9��9S��9���9?��9Ҷ�9@��9��9���9���9~��9���9
��9޲�9���9T��9���9%��9e��9x   x   ���9��9G��97��9��9���9���9%��9w��9���9z��9ô�9��9B��9���9��9��9R��9��9���9���9���9���9���9���9p��9���9��9��9��9x   x   Y��9ֳ�9x��9ϵ�9Ѵ�9��9h��9δ�9���9���9���9��9"��9���9=��9���9���9���9���9 ��9���9��9���9#��9/��9/��99��9���9���9δ�9x   x   ��9��9̲�9���9���9���9���9��9ʷ�9*��9���9ҳ�9���9Ƴ�9��9��9K��9.��9��9���9��9ݲ�9���93��9���9(��9���9���9Z��9���9x   x   ,��9Ҹ�9���9���9���9��99��9��9y��9��9���94��9u��9���9Ӳ�9ݵ�9X��9.��9/��9\��9���9���9p��9,��9(��9з�9 ��9��9��9E��9x   x   ɮ�9!��9��9;��9'��9ذ�9(��9���9���9��9V��91��9
��9m��9���9���9���9+��9���9Y��9i��9Y��9���93��9���9��9ư�9ر�9��9��9x   x   ���9��9���9��9���9|��9˷�9Q��9���9#��9յ�9���9m��9���9��9��9���9��9e��9���9���9���9��9���9���9޲�9ر�9W��93��9x��9x   x   ���9���9=��9-��9i��9���9=��9���9��9Է�9G��9V��91��9���9s��9��9���9���9ִ�9��9���9#��9��9���9\��9��9��99��9���9���9x   x   ���9̲�9���9`��9ٲ�9���9Q��9>��9���9��9Y��9��9���9��9��9���9³�9Z��9ٲ�9���9'��9h��9��9δ�9���9D��9��9|��9���9,��9x   x   ���9��9��9���9��9f��9���9��9]��9���9��9���9���9k��9!��9���9���9���9&��9���9T��9d��9���9��9��9���9���9���9��9��9x   x   ��9k��95��9!��9P��9p��9���9��9���9��9��9��9���9P��9G��9���9L��9��9F��9���9���9���9���9���9���9���9���9��9���9���9x   x   ��92��9���9���9��9@��9o��9���9���9���9g��9Z��9���9b��9=��9+��9���9��9���9���9O��9���9���9��9��9���9���9���9��9	��9x   x   ���9��9���9g��9^��9���9w��9.��9*��9v��9���9���9���9>��9���9���9���9���9k��9���9H��9���95��9#��9���9j��9<��9���9+��9K��9x   x   ��9R��9��9d��9���9���9���9s��9��9���9���9<��9��9��9:��9���9���9f��9���9���94��9���9H��9-��9���9���9���9��9��9k��9x   x   g��9l��9B��9���9���9)��9��9z��9���9���9��9���9H��9��9���9��9���9���9���9u��9���9���9���91��9���9���9H��9���9���9���9x   x   ���9���9p��9u��9���9��9h��9���9��9b��9���9���9m��9���9��9���9���9���9)��9���9���9��9���9<��9��9���9a��9H��9F��9.��9x   x   
��9��9���9,��9t��9x��9���9\��9���9U��9���9C��9���9���9<��9*��9y��9���9���9G��9���9��9g��9d��9k��9��9��9���9���9s��9x   x   Z��9���9���9)��9��9���9��9���9L��96��9��9,��9B��9��9���9���9���9(��9P��9���9���9��9���9<��9}��9���9���92��9��9���9x   x   ���9��9���9r��9���9���9a��9S��95��9���9���9���9���9\��9E��9���9���9*��9���9��9���9���94��9���9���9���9l��9���9���9���9x   x   ��9���9i��9���9��9��9���9���9��9���9���9\��9��9���9��9&��9M��9��97��9���9���9��9[��9q��9��9V��9���9h��9%��9b��9x   x   ���9	��9Y��9���9<��9���9���9>��9&��9���9X��9���9y��9_��9���9��9��9���9���9���9"��9���9���9���9��9���9���9���9���9&��9x   x   ���9���9���9���9��9F��9t��9���9D��9���9��9~��9���94��9���9��9��9���9���9���9o��90��9���93��9���9T��9T��9p��9��9��9x   x   k��9T��9e��9B��9��9��9���9���9��9W��9���9^��97��9���9{��9l��9���9Q��9^��9Z��9��9Y��9��9P��9���9���9��9���9$��9���9x   x   ��9D��9:��9���9;��9���9��9:��9���9G��9��9���9���9z��9���9}��9��9���9O��9m��9���9O��9���9��9H��9]��9���9���9n��9���9x   x   ���9���9.��9���9���9	��9���9/��9���9���9*��9��9y��9i��9���9���9b��9���9_��9D��9���9��9^��9*��9���9���9���9��9���9���9x   x   ���9N��9���9���9���9���9���9x��9���9���9K��9 ��9��9���9!��9d��9]��9���9���9���9X��9,��9���9���9��9���9:��9���9#��9A��9x   x   ���9��9��9���9f��9���9���9���9+��9.��9��9���9���9R��9���9���9���9���9���9���9S��9z��9���9���9���9���9���9���9���9d��9x   x   %��9D��9���9e��9���9���9(��9���9J��9���98��9���9���9_��9L��9`��9���9���9!��9��9���9���9���9���9���9���9���9o��9��9���9x   x   ���9���9���9���9���9n��9���9F��9���9��9���9���9���9W��9j��9D��9���9���9��9���9���9N��9��9;��9��9���9���9���9���9���9x   x   V��9���9M��9H��94��9}��9���9���9���9���9���9"��9n��9��9��9���9Z��9R��9���9���9Q��9W��9\��9s��9���9���9���9���9���9s��9x   x   c��9��9���9���9���9���9��9��9��9���9��9~��9/��9X��9N��9��9'��9{��9��9N��9V��9f��9���9A��9Q��9
��9$��9��9���9���9x   x   ���9���9���9;��9G��9���9���9j��9���94��9\��9���9���9
��9���9^��9���9���9���9��9\��9���9���9#��9e��9}��9���9���9���9���9x   x   ��9���9
��9#��9*��90��9:��9a��9;��9���9o��9���93��9Q��9��9)��9���9���9���9;��9u��9E��9 ��9R��9���9���9?��9���9���9���9x   x   ���9���9��9���9���9���9��9p��9|��9���9��9��9���9���9G��9���9��9���9���9��9���9S��9`��9���9"��9���9���9v��9��9���9x   x   ���9���9���9k��9���9���9���9��9���9���9V��9���9U��9���9]��9���9���9���9���9���9���9��9z��9���9���9}��9���9^��9���9m��9x   x   ���9���9���9=��9���9G��9b��9	��9���9l��9���9���9Q��9	��9���9���9:��9���9���9���9���9$��9���9>��9���9���9���9B��9���9��9x   x   ���9��9���9���9 ��9���9K��9���93��9���9i��9���9p��9���9���9��9���9���9q��9���9���9��9���9���9y��9c��9A��9F��9���9"��9x   x   ��9���9��9+��9��9���9F��9���9��9���9"��9���9��9��9o��9���9"��9���9��9���9���9���9���9���9��9���9���9���91��9���9x   x   ��9���9��9L��9o��9���9.��9s��9���9���9c��9(��9
��9���9���9���9A��9d��9���9���9u��9���9���9���9���9r��9"��9!��9���9���9x   x   ���9B��9���9,��9
��9`��9`��9i��96��9���9Y��9���9d��9���9��9+��9���9���9���9���9���9���9���9���9��9���9���9���9n��9F��9x   x   D��9"��9���9H��9K��9��9���9���9���9���9��9���9���9g��9���9���9���9G��9���9��9d��9@��9���9���9t��9J��9���9���99��9���9x   x   ���9���9A��9��9���9���9K��9��9���9���9t��9%��9���9��9���9���9y��9*��9���9���9���9D��93��9���9Z��9���9���9���9��9y��9x   x   -��9K��9��9��9m��9`��9:��93��9G��9���9���9���9���9"��9���9,��9!��95��9"��9W��9#��9z��9b��9.��9���9P��9���9���9)��9Q��9x   x   ��9I��9���9j��9���9���9���9���9���9���9���9���9���9���9��91��9���9���9.��9���9���9���9��9$��9��9���9e��9��9��9���9x   x   a��9	��9���9^��9���9���9��9���9���9��9���9s��9��9Z��94��9"��9	��9���9���9���9z��9���9���9���9��9^��9���9u��9���9���9x   x   b��9���9L��9<��9���9��9a��9���9���9z��9F��9���9���9>��9f��9���9F��9h��9���9���9@��9���9���9��9���9��9���9e��9���9��9x   x   h��9���9��95��9���9���9���9��9���9|��9���9���9���9	��9u��9#��9��9���9q��9���9���9;��9B��9���9��9%��9���9��9F��9&��9x   x   8��9���9���9H��9���9���9���9���9���9���9���9���9 ��9i��9��9a��9���95��9���9��9	��9k��9n��9]��9��9"��9 ��9��9���9���9x   x   ���9���9���9���9���9!��9w��9|��9���9Z��9j��9���9Z��9���9X��9C��9���9H��9���9W��9A��9���9���9U��9
��9n��9)��9��9���9���9x   x   ]��9��9u��9���9���9���9G��9���9���9p��9 ��9>��9���9���9}��9���9B��9M��9��9|��9��9)��97��9���9C��9���9��9n��9���9��9x   x   ���9���9$��9���9���9u��9���9���9���9���96��9{��9���9���9���9��9O��9���9V��9���9���9z��9���9���9���9���9|��9���9���9E��9x   x   d��9���9���9���9���9��9���9���9��9[��9���9���9���90��9��9���96��9r��9���9%��9x��9���9v��9���9���9���9��9���9���9���9x   x   ���9h��9��9��9���9\��9>��9��9i��9���9���9���91��9���9��9���9���9'��9���9O��9���9Q��9^��9���9&��9���9<��9>��9	��9���9x   x   ��9���9���9���9��98��9c��9s��9��9V��9{��9���9��9��9���9 ��9���9���9��96��9���9���9.��9���9r��9���9B��9���9���9v��9x   x   .��9���9���9-��9.��9"��9���9%��9c��9D��9���9!��9���9���9$��9:��9o��9���9���9:��9(��9���9���9Q��9 ��9���9��9j��9���9��9x   x   ���9���9v��9$��9���9��9?��9��9���9���9@��9S��96��9���9���9k��9���9a��9���9��9P��9���9���9���9���9`��9S��9^��9���9$��9x   x   ���9K��9)��9:��9���9���9g��9���93��9K��9R��9���9v��9%��9���9���9_��9���9&��9i��9>��9~��9���9���9���9���9���9D��9��9��9x   x   ���9���9���9!��9-��9���9���9q��9���9���9��9U��9���9���9��9���9���9(��9��9<��9���9M��9w��9���9���9)��9o��95��9	��9��9x   x   ���9��9���9Z��9���9���9���9���9��9T��9}��9���9'��9O��94��99��9��9h��9<��9���9��9d��9���9���9���9���9���9,��9k��9��9x   x   ���9_��9���9%��9���9~��9A��9���9��9A��9��9���9{��9���9���9&��9N��9=��9���9��9���9���9F��9E��9E��9���9���99��9���9|��9x   x   ���9@��9D��9{��9���9���9���98��9k��9���9*��9{��9���9Q��9���9���9���9~��9N��9e��9���9?��9��9���9���9:��9���9��9���9���9x   x   ���9���90��9a��9��9���9���9B��9n��9���96��9���9u��9Z��9-��9���9���9���9x��9���9G��9��9���9n��9`��9���9���9���9���9���9x   x   ���9���9���9+��9'��9���9 ��9���9]��9T��9��9���9���9���9���9R��9���9���9���9���9C��9���9m��96��9���9+��9���9���9���9V��9x   x   ~��9u��9\��9���9��9��9���9��9��9
��9F��9���9���9'��9s��9��9���9���9���9���9F��9���9b��9���9���9��9w��9L��9l��9��9x   x   ���9H��9���9M��9���9_��9
��9%��9$��9m��9���9���9���9���9���9���9`��9���9'��9���9���99��9���9,��9��9*��9��9h��9���9}��9x   x   ���9���9���9���9e��9���9���9���9 ��9&��9��9}��9��9:��9?��9��9S��9���9j��9���9���9���9���9���9s��9��9���9���9���91��9x   x   ���9���9���9���9��9q��9g��9��9��9���9m��9���9���9B��9���9i��9Z��9E��93��9-��9>��9��9���9���9I��9e��9���9���9���9g��9x   x   l��9:��9��9)��9 ��9���9���9E��9���9���9���9���9���9��9 ��9���9���9��9��9j��9���9���9���9���9l��9���9���9���9X��9t��9x   x   C��9���9t��9R��9���9���9 ��9&��9���9���9��9F��9���9���9t��9���9%��9��9��9��9{��9���9���9U��9��9{��94��9g��9s��9o��9x   x   ��9��9��9v�9X�9�9�
�9v�9~�9�	�9�	�9��9��9��9i
�9��9��9U�9u�9��9"	�9�
�9�9�
�9��9��9��9I�9	�9	�9x   x   ��9�
�9��9W	�9m
�9;�9��9r
�9Y�9��9�
�9��9�
�9�9��9��9,
�9�
�9d�9o
�9c�9�
�9p�9��9v�9�	�9�	�9��9F
�9�	�9x   x   ��9��9�
�9m�9W�9�	�9
�9u	�9t�9�
�9P�9b�90	�9��9s�9��9
�9R�9 �9]�9-�9X�92	�9}
�9F�96�9:�9"�9��9R	�9x   x   x�9W	�9m�9�
�9��9�9-�9D�9�9*�9�
�9�
�9��9�	�9��9P�9b	�9��9�9�	�9Z�9��9H�9��9�
�9��9��9��9��9��9x   x   X�9i
�9U�9��9T�9�
�9��9%�9�	�9�
�9�
�9r
�9�9=�9��9T�9�9�	�9w�9�
�9�
�9=�9��9��9��9�
�9��9��9��9��9x   x   �9=�9 
�9�9�
�9e�94
�9j�9w
�9��9d�9��9�9��9��9��9 �9�	�9��9�
�9G�9�	�9��9v	�9��9#�9z�9��9��9m�9x   x   �
�9��9
�9/�9��9:
�95�9��9��9��9_�9��9c	�9��9��9*�9��9��9-�9
�9��9J�9�	�9`�9�
�9�9��9��92�9��9x   x   v�9q
�9t	�9E�9�9n�9��9��9��9H
�9��9M�92�9��9?
�9\�9��9y�9��9y
�9��9u	�9�
�9	�9��9�
�9Q�9�9�
�9��9x   x   ~�9Z�9t�9�9�	�9v
�9��9��9V	�9>�9��9 �9|�94�9u
�9�9��99
�9I�9 �9��9a�9�9�
�9�
�9��9��9��9 �9
�9x   x   �	�9��9�
�9)�9�
�9��9��9K
�98�9��9��9��9j�9h�9��9��9��9�	�9
�95�9g�9"
�9��9t�9�
�9�
�9M�9^
�9��9��9x   x   �	�9�
�9P�9�
�9�
�9e�9^�9��9��9��9��9p�9��9��91�9y�9��9��9��9�	�9�	�9�	�9V�9��9e�9��9r�9��9C�9[	�9x   x   ��9��9`�9�
�9r
�9��9��9T�9��9��9u�9\�9y�9�9��9�
�9J	�9�
�9}�9��9[�9 �9�
�9q
�9?
�9�	�9�
�9|
�9Q�9��9x   x   ��9�
�9-	�9��9�9�9`	�92�9s�9i�9��9q�9F	�9��9z�9��9�
�9�
�9��9��9/�9��9��9m
�9�9�
�9,�9!	�9n
�92�9x   x   ��9�9��9�	�9=�9��9��9��92�9l�9��9�9��9o�9r	�9q�9�
�9��9>
�9$
�9�
�9��9��9S�9[�9_�90	�9�
�9�	�9S
�9x   x   d
�9��9y�9��9��9��9��9B
�9s
�9��96�9��9w�9p	�9 	�9��9O�9��9$�9F�9b�9Q
�9�9��9��9�
�9��9*�9�
�9��9x   x   ��9��9��9Q�9R�9��9*�9Y�9	�9��9y�9�
�9��9l�9��9��9/�9@	�9��9�9��9#�9�9T�9'�99�9��9�9n	�9F�9x   x   ��9,
�9
�9e	�9
�9$�9��9��9��9��9��9H	�9�
�9�
�9T�92�9G
�9�	�9�
�9�
�9��9"
�9�9�	�9�9J�9�
�9V
�9��9�
�9x   x   U�9�
�9L�9��9�	�9�	�9��9x�97
�9�	�9��9�
�9�
�9��9��9?	�9�	�9-�9r�9�
�9��9��9��9��9,
�9C�9��9
�9�
�9��9x   x   s�9f�9��9�9x�9��9*�9��9J�9
�9��9|�9��99
�9 �9��9�
�9r�9�	�9��9�	�9��9��9!�9L
�91�9v
�9n�9�
�9
�9x   x   ��9o
�9^�9�	�9�
�9�
�9�	�9x
�9 �95�9�	�9��9��9&
�9I�9�9�
�9�
�9��99	�9��9�	�99	�9��9�	�9�
�99�9w�9�
�9��9x   x   $	�9d�91�9U�9�
�9G�9��9��9��9h�9�	�9Z�9*�9�
�9b�9��9��9��9�	�9��9�
�9��9�	�9p�9s	�9��9��9B
�9<
�9��9x   x   �
�9�
�9]�9��9<�9�	�9L�9y	�9_�9#
�9�	�9�9��9��9S
�9$�9$
�9��9��9�	�9��93�9��9%	�9r�9�
�9/	�9�	�9C�9�	�9x   x   �9l�91	�9G�9��9��9�	�9�
�9�9��9S�9�
�9��9��9�9�9�9��9��99	�9�	�9��9	�9�9��9.�9��9�
�9��9|�9x   x   �
�9��9}
�9��9��9u	�9e�9�9�
�9t�9��9s
�9q
�9V�9��9T�9�	�9��9�9��9r�9&	�9�9�9a�9v�9�
�9+	�9��9�
�9x   x   ��9p�9G�9�
�9��9��9�
�9��9�
�9�
�9a�9;
�9�9\�9��9&�9��90
�9N
�9�	�9p	�9p�9��9_�9P�9�	�9�9H
�9<
�9�	�9x   x   ��9�	�97�9��9�
�9%�9�9�
�9��9�
�9��9�	�9�
�9_�9�
�95�9J�9?�9/�9�
�9��9�
�9-�9q�9�	�9�9�9�	�9
�9�
�9x   x   ��9�	�97�9��9��9|�9��9I�9��9O�9s�9�
�9.�95	�9��9��9�
�9��9v
�9:�9��90	�9��9�
�9�9�9�9W�9m�9�9x   x   H�9��9 �9��9��9��9��9��9��9^
�9��9{
�9	�9�
�9.�9�9S
�9
�9r�9x�9B
�9�	�9�
�9,	�9G
�9�	�9Y�9��9��9o�9x   x   	�9H
�9��9}�9��9��92�9�
�9!�9��9B�9Q�9j
�9�	�9�
�9q	�9��9�
�9�
�9 �9=
�9D�9��9��9=
�9
�9q�9��9s�9��9x   x   	�9�	�9W	�9��9��9l�9��9��9
�9��9Y	�9��91�9O
�9��9K�9�
�9��9
�9��9��9�	�9z�9�
�9�	�9�
�9�9r�9~�9��9x   x   '(�9�,�9*�9�*�9.�9Y(�9*�9-�9�(�9�+�9�)�9N&�9�*�9u)�9�(�9�,�9�)�9�)�9�*�9'�9e)�9q-�9>(�9l+�9(*�9�'�9E/�9�*�9�+�9�,�9x   x   �,�9F.�9i&�9e,�9�*�9�(�93-�9�+�9J)�9�(�9!*�9S*�9*�9p,�9)*�9�*�9+�9*�9k*�93*�9�'�9�(�9�-�9M-�9Y)�9�)�9,�9H%�9m-�9�-�9x   x   *�9k&�9g+�9�-�9�+�9I-�9|,�9*�9�+�9�)�9w,�9�*�9�+�9�+�9�*�9�+�9-�9�*�9�+�9�*�9P,�91)�9�+�9�,�9T,�9 .�9�,�94'�9b)�9�&�9x   x   �*�9c,�9�-�9P)�9#,�9�(�9�$�9�*�9>)�9+�9*�98,�9<*�9�+�9�+�9*�9�*�9J+�9|*�9�'�9�+�9�$�9/*�9E+�9�)�9-�9+�9�+�9�(�9�(�9x   x   .�9�*�9�+�9$,�9�-�9*�9�+�9�(�9',�9�+�9-'�9�(�9�'�9�*�9 (�9)�9�'�9_+�9�-�9(�9�+�9�)�9�-�9�,�9�+�9/,�9�-�9�-�94)�91.�9x   x   Y(�9�(�9K-�9�(�9!*�9�2�9�(�9+�9+�9>*�9�.�9�,�9�*�9k*�9G,�9�/�9l)�9*�94+�9�(�9Y3�9�)�9;)�9�,�9(�9(�9�.�9N)�9�(�9u.�9x   x   *�93-�9z,�9�$�9�+�9�(�9(�9/�9�'�9�-�9�-�9u+�9o+�9�+�9�-�9<-�9�)�9�.�9M(�9�'�9E,�9%�9�+�9�.�9�)�9W*�9�)�9�#�9�*�9�)�9x   x   -�9�+�9*�9�*�9�(�9+�9/�9m/�9�*�9�*�9�)�9^(�9V(�9�)�9�*�9�)�9�.�9=/�9�+�9�(�9�)�9L*�9<+�9b,�9q-�9�*�9*�9T)�9�*�9;-�9x   x   �(�9K)�9�+�9B)�9+,�9+�9�'�9�*�9)(�9,�9�)�9�&�9\)�9�+�9h)�9�*�9�(�9$*�9O,�9�)�9�+�9�)�9�(�9V*�9�*�9�)�9�2�9�)�9�+�9�)�9x   x   �+�9�(�9�)�9+�9�+�9>*�9�-�9}*�9,�9N+�9r+�9G+�9�+�9f+�9�)�9t-�90*�9�+�9�)�9�)�9�'�9,�9�(�9c)�9W+�9�+�9�,�9d*�9�)�9)�9x   x   �)�9&*�9z,�9*�9('�9�.�9�-�9�)�9�)�9q+�9�2�9m+�9�)�9�)�9F.�96.�9M'�9'+�9�,�9�)�9�*�90�9�'�9�+�9�*�9Q&�96*�9L,�9(�9�/�9x   x   J&�9T*�9�*�98,�9�(�9�,�9t+�9](�9�&�9K+�9o+�9�%�9�(�9�*�9:-�9�)�9t*�9(*�9#*�9�&�9�(�9-)�9,�9 ,�9{-�9@-�9	-�9 +�9�(�9�)�9x   x   �*�9*�9�+�9:*�9�'�9�*�9q+�9T(�9^)�9�+�9�)�9�(�9�+�9�*�9\&�9�*�9*-�9}*�9�*�9�)�9+�9�*�9�*�97*�9�1�9�)�9:*�9�,�9)*�9*�9x   x   q)�9v,�9�+�9�+�9�*�9p*�9�+�9�)�9�+�9a+�9�)�9�*�9�*�9�+�9�+�9�*�95+�9%)�9)�9.+�9�,�9�,�9S)�9-)�9�)�9�)�9",�9�+�9:+�9+)�9x   x   �(�9'*�9�*�9~+�9#(�9J,�9�-�9�*�9j)�9�)�9E.�97-�9a&�9�+�9�+�9�*�9�)�9�)�9�,�9�)�9C'�9�,�9�*�9(�9�)�9�,�9'�9]+�9A,�9')�9x   x   �,�9�*�9�+�9*�9)�9�/�98-�9�)�9�*�9p-�93.�9�)�9�*�9�*�9�*�9�+�9�+�9#+�9�-�9�*�9�)�9�+�9*�9�*�9�+�9:*�9x)�9�,�9�,�9�,�9x   x   �)�9+�9-�9�*�9'�9l)�9�)�9�.�9�(�92*�9N'�9u*�9.-�95+�9�)�9�+�9�-�95,�9�)�9�,�9O+�9�+�9f'�9M,�9p*�97-�9]+�9�,�9<+�9�*�9x   x   �)�9*�9�*�9J+�9[+�9*�9�.�97/�9 *�9�+�9(+�9+*�9z*�9$)�9�)�9'+�9<,�9�&�9*�9�+�9�*�9s+�94*�9�*�9F+�9)�9 &�9�,�9�-�9Y)�9x   x   �*�9m*�9�+�9*�9�-�94+�9R(�9�+�9M,�9�)�9�,�9"*�9�*�9)�9�,�9�-�9�)�9 *�9,-�9�(�9�*�9.�9�*�9)�9�-�9P*�95*�9n,�9L+�9�)�9x   x   '�93*�9�*�9�'�9(�9�(�9�'�9�(�9�)�9�)�9�)�9�&�9�)�93+�9�)�9�*�9�,�9�+�9�(�9/.�9x.�9G/�9�,�9�'�9�+�9|,�9)+�9�*�9M,�9�(�9x   x   c)�9�'�9O,�9�+�9�+�9[3�9I,�9�)�9�+�9�'�9�*�9�(�9+�9�,�9A'�9�)�9N+�9�*�9�*�9x.�9�&�9�.�9�,�9v*�90+�9)�9�&�9l+�9�*�9�)�9x   x   q-�9�(�90)�9�$�9�)�9�)�9#%�9L*�9�)�9,�90�92)�9�*�9�,�9�,�9�+�9�+�9u+�9!.�9F/�9�.�9�,�9\*�9�+�9f,�9,-�9�,�9,,�9*)�9�/�9x   x   ;(�9�-�9�+�9/*�9�-�99)�9�+�97+�9�(�9�(�9�'�9	,�9�*�9S)�9�*�9*�9h'�95*�9�*�9�,�9�,�9X*�9�(�9�)�9�)�9`)�9�*�9+�9�'�9�(�9x   x   m+�9P-�9�,�9D+�9�,�9�,�9�.�9`,�9U*�9e)�9�+�9�+�93*�9+)�9(�9�*�9M,�9�*�9)�9�'�9y*�9�+�9�)�9s)�9G)�9Q*�9:,�9-�9�)�9�*�9x   x   &*�9Y)�9X,�9�)�9�+�9(�9�)�9r-�9�*�9U+�9�*�9-�9�1�9�)�9�)�9�+�9o*�9H+�9�-�9�+�9/+�9j,�9�)�9J)�9{1�9_-�9*�9	*�9s*�9�.�9x   x   �'�9�)�9�-�9-�9/,�9(�9U*�9�*�9�)�9�+�9T&�9D-�9�)�9�)�9�,�9;*�95-�9)�9R*�9|,�9)�9.-�9_)�9V*�9`-�9�&�9T,�9�+�9�)�9�)�9x   x   F/�9,�9�,�9+�9�-�9�.�9�)�9
*�9�2�9�,�96*�9-�96*�9#,�9'�9z)�9^+�9&�94*�9*+�9�&�9�,�9�*�9;,�9*�9S,�921�9�)�9=+�9r.�9x   x   �*�9J%�97'�9�+�9�-�9L)�9�#�9[)�9�)�9e*�9M,�9�*�9�,�9�+�9Z+�9�,�9�,�9�,�9l,�9�*�9f+�9-,�9+�9-�9
*�9�+�9�)�9�"�9�(�9-�9x   x   �+�9g-�9^)�9�(�91)�9�(�9�*�9�*�9�+�9�)�9(�9�(�9+*�9>+�9D,�9�,�9;+�9�-�9R+�9O,�9�*�9,)�9�'�9�)�9r*�9�)�9;+�9�(�9�*�9T(�9x   x   �,�9�-�9�&�9�(�92.�9w.�9�)�9;-�9�)�9)�9�/�9�)�9*�9/)�9%)�9�,�9�*�9[)�9�)�9�(�9�)�9�/�9�(�9�*�9�.�9�)�9w.�9-�9R(�9�%�9x   x   �F�9K�9�K�9KI�9�H�9RK�9N�9�G�9L�9�J�9PM�9�L�9�K�9-M�90L�9&K�9L�9�L�9dL�9FM�9�L�9�L�9K�9�F�9�M�9�I�9XJ�9�I�9�L�9-K�9x   x   K�9J�9M�9�K�9J�9WL�9�J�9�I�9�M�9�L�9�P�92L�9L�9yL�9�J�9�K�9kL�9�K�9�K�9�P�9L�9_M�9�J�9~J�9�M�9(J�9�J�9eL�9GI�9�K�9x   x   �K�9M�9L�9@J�9�I�9�H�9UN�9�M�9�J�9.L�9�H�90J�9�I�9I�9+M�9BH�9qJ�9,J�9�H�9:M�9�J�9qM�9�M�9�G�9�I�9nJ�9YM�9�M�9LK�9�P�9x   x   LI�9�K�9?J�9J�9�J�9�K�9kO�9�J�90M�9�K�9L�9�O�9�H�9PM�9�M�9MI�9O�9�L�9�J�9�L�9�K�9O�9�M�9uJ�9pJ�9�I�9�I�9J�9�L�9�L�9x   x   �H�9~J�9�I�9�J�9L�9]J�9mK�9UM�9�J�9M�93M�9�N�9�M�9�J�9�M�9uN�90M�9iM�9+L�9�L�9�K�96I�9~K�9�K�91I�9}L�9%I�9�K�9�L�9�L�9x   x   RK�9UL�9�H�9�K�9]J�9H�9�M�9�I�9�J�9L�9�D�9FL�9�H�9qH�9L�9bE�9`K�9%J�9�I�9�M�9jI�9�J�9�K�9�H�9�K�9(J�9�I�9�N�9�M�9�I�9x   x   N�9�J�9XN�9lO�9nK�9�M�9kL�9�I�9
N�9.L�9�J�9IM�9YM�9�M�9wJ�9L�9FO�9#I�9jM�9~L�9�J�9�O�9xM�9�K�9 N�9cI�9hK�9O�9rL�9�H�9x   x   �G�9�I�9�M�9�J�9TM�9�I�9�I�9�F�9#I�9eM�9�G�90N�9�M�9�G�9�M�9vH�9�F�97I�9tJ�9;N�9�I�9�N�9�H�9�F�9K�9M�9BL�9�K�91M�9�J�9x   x   L�9�M�9�J�90M�9�J�9�J�9N�9#I�9sN�9�J�9.K�9R�9xK�9�J�9�N�9�H�9O�9�I�9�J�9�M�9_J�9:N�9�L�9�L�9�K�9J�9~G�9wI�9�L�9�L�9x   x   �J�9�L�9+L�9�K�9M�9L�9,L�9dM�9�J�96N�9L�9�K�9
N�9�I�9�M�9dK�9�L�9cN�9�J�9�L�9�K�9�J�9L�9;M�9M�9I�9�J�9zL�9�L�9UL�9x   x   NM�9�P�9�H�9	L�93M�9�D�9�J�9�G�9.K�9L�9�@�9L�9L�9�G�9PK�9RD�9	L�9�L�9�H�9�P�9/N�9%K�9�J�9L�9�L�9L�9�K�9�L�9QK�9IK�9x   x   �L�9.L�90J�9�O�9�N�9CL�9JM�9)N�9R�9�K�9L�9Q�9N�9�L�9�L�9�O�9�N�9�J�9=K�9]L�9?J�9^L�9"N�9I�9^I�9�I�9/J�9�L�9oK�9�J�9x   x   �K�9L�9�I�9�H�9�M�9�H�9[M�9�M�9{K�9N�9L�9N�9$N�9PH�9�K�9�I�9�I�9xL�9M�9yM�9�L�9�J�9�I�9nJ�9�I�9�I�9I�9HM�9�L�9=M�9x   x   *M�9wL�9I�9TM�9�J�9jH�9�M�9�G�9�J�9�I�9�G�9�L�9OH�9M�9EM�9�H�9!L�9+L�9#M�9?J�9M�91L�9EL�9nM�9�M�9%M�9HK�9FK�9�J�9N�9x   x   -L�9�J�90M�9�M�9�M�9L�9yJ�9�M�9�N�9�M�9RK�9�L�9�K�9FM�9�L�9pK�9�L�9�M�9�K�9�H�9�L�9CL�9nJ�9�M�9�I�9�L�9�M�9�J�9yJ�9M�9x   x   'K�9�K�9BH�9NI�9vN�9cE�9L�9xH�9I�9fK�9VD�9�O�9�I�9�H�9rK�9�I�9�J�9�G�9�K�9�L�9�K�9�I�9oN�9�N�9I�9�K�9nK�9�J�9J�9�J�9x   x   L�9iL�9oJ�9O�9/M�9^K�9DO�9�F�9O�9�L�9L�9�N�9�I�9 L�9�L�9�J�9�J�9�K�9�K�9�K�9L�9NM�9wK�9lN�9 L�9+L�9�L�9�K�9�H�9UJ�9x   x   �L�9�K�9,J�9�L�9mM�9*J�9'I�9;I�9�I�9eN�9�L�9J�9wL�9*L�9�M�9�G�9�K�9N�9�K�9�J�9�L�9eL�9|J�9:L�9ZJ�9K�9XM�9 L�9]J�9�M�9x   x   fL�9�K�9�H�9�J�9)L�9�I�9lM�9rJ�9�J�9~J�9�H�9=K�9M�9!M�9�K�9�K�9�K�9�K�9vL�9L�9�H�9J�9�J�9�L�9�L�9dK�9�L�9*J�9J�9�M�9x   x   FM�9�P�9:M�9�L�9�L�9�M�9yL�99N�9�M�9�L�9�P�9YL�9vM�9=J�9�H�9�L�9�K�9�J�9L�9�L�9�I�9rI�9K�9_K�91K�9K�9�L�9�J�9OK�9XL�9x   x   �L�9L�9�J�9�K�9�K�9jI�9�J�9�I�9`J�9�K�94N�9>J�9�L�9M�9�L�9�K�9L�9�L�9�H�9�I�9tH�9�I�9wK�9SL�9;L�9�K�9�L�9�K�9xL�9ZK�9x   x   �L�9`M�9qM�9�N�90I�9�J�9�O�9�N�9<N�9�J�9#K�9^L�9�J�91L�9AL�9�I�9PM�9dL�9J�9pI�9�I�9�H�9�J�9vM�9�I�9mL�9>L�9HL�9(L�9|J�9x   x   K�9�J�9�M�9�M�9�K�9�K�9wM�9�H�9�L�9L�9�J�9N�9�I�9FL�9mJ�9pN�9vK�9{J�9�J�9K�9vK�9�J�9,M�9�M�9J�9|L�9dI�9�L�9CK�9�K�9x   x   �F�9|J�9�G�9sJ�9�K�9�H�9�K�9�F�9�L�9<M�9L�9I�9oJ�9jM�9�M�9�N�9jN�97L�9�L�9\K�9TL�9tM�9�M�9�N�9M�9{J�9�I�9M�9	M�9�M�9x   x   �M�9�M�9�I�9rJ�90I�9�K�9!N�9K�9�K�9M�9�L�9\I�9�I�9�M�9�I�9	I�9#L�9ZJ�9�L�9-K�99L�9�I�9J�9M�9J�9+I�9[L�9�K�9�K�9�K�9x   x   �I�9&J�9oJ�9�I�9~L�9*J�9`I�9M�9J�9 I�9L�9�I�9�I�9$M�9�L�9�K�9+L�9K�9eK�9K�9�K�9jL�9{L�9{J�9)I�9SL�9J�9�K�9�K�9�I�9x   x   [J�9�J�9WM�9�I�9%I�9�I�9hK�9AL�9|G�9�J�9�K�90J�9
I�9HK�9�M�9mK�9�L�9XM�9�L�9�L�9�L�9>L�9aI�9�I�9ZL�9J�9�E�9ML�9�L�9�I�9x   x   �I�9gL�9�M�9J�9�K�9�N�9O�9�K�9uI�9{L�9�L�9�L�9JM�9GK�9�J�9�J�9�K�9L�9+J�9�J�9�K�9JL�9�L�9M�9�K�9�K�9KL�9�N�9�M�9K�9x   x   �L�9FI�9KK�9�L�9�L�9�M�9pL�93M�9�L�9�L�9QK�9kK�9�L�9�J�9wJ�9J�9�H�9`J�9J�9QK�9vL�9'L�9EK�9
M�9�K�9�K�9�L�9�M�9EN�99L�9x   x   0K�9�K�9�P�9�L�9�L�9�I�9�H�9�J�9�L�9RL�9IK�9�J�9=M�9N�9M�9�J�9YJ�9�M�9�M�9[L�9WK�9|J�9�K�9�M�9�K�9�I�9�I�9K�9<L�9zP�9x   x   It�9�l�9m�9�n�9wm�9�r�9�o�91o�9�q�9'j�9ml�9�m�9�k�9xk�9�n�9)n�9�m�9kk�9�l�9�m�9Vl�9�j�9�p�9�o�9�n�9�p�9\o�9�o�9�l�9�l�9x   x   �l�9Lk�9{q�9�n�9o�9�m�9�m�9m�9�o�9l�9yj�9�n�9�n�9mm�9�n�9o�9an�9�n�9�m�9Qj�9l�9�o�9�m�9�m�9�o�9;o�9m�9Tq�96k�9wm�9x   x   m�9{q�9i�9:m�9�q�9�m�9�j�9<j�9m�9Hm�9�m�9�o�9�o�9�q�9m�9�p�9o�97p�9�n�9]m�9�l�9�j�9Wj�9m�9�p�9[m�9fj�9r�9l�9Qk�9x   x   �n�9�n�9<m�9�p�9o�9�l�9�o�9*l�9So�9�n�9Om�90i�9�m�9$k�9�k�9�n�9wi�9�l�9�m�9�o�9Rl�9�o�9gn�9�n�9dq�9m�9�l�9�o�9�m�9/m�9x   x   wm�9o�9�q�9o�9Ll�9�p�9%m�9�n�9�k�9�k�9�n�9cn�9p�9o�9xo�94n�9�n�9l�9Cl�9an�9|m�9�o�9�k�9ao�95p�9�p�9qn�9=k�9�j�9�l�9x   x   �r�9�m�9�m�9�l�9�p�9'i�9�m�9Ro�9�m�9=o�9=n�9Yl�9�p�9�p�9l�9Qn�9So�9�m�9$o�9xm�9�i�9^q�9�l�9�n�9�m�9'q�9n�9�k�9�j�9�m�9x   x   �o�9�m�9�j�9�o�9!m�9�m�9p�9�m�9�p�9l�9�n�9�l�9�k�9Jm�9�n�9�k�9�p�93m�9�p�9m�9�l�9
p�9�i�9�n�9�o�9p�9Pl�9�o�9�l�9o�9x   x   /o�9m�9<j�9)l�9�n�9Uo�9�m�9 p�9!o�9im�9)r�9�k�9k�9uq�9n�9.o�9�p�9Km�9ao�9jo�9�k�99k�9�l�9�n�9�k�9�n�9n�9n�9�o�9�k�9x   x   �q�9�o�9m�9To�9�k�9�m�9�p�9'o�9eo�9=m�9�m�9Lj�9�n�9cm�9�n�9�n�9q�95m�9�k�9�o�9Ol�9p�9)r�9�n�9ej�9)q�9Xm�9�o�9k�9.o�9x   x   +j�9l�9Pm�9�n�9�k�9>o�9l�9jm�98m�9rl�9�m�9$m�9�k�9m�9xn�9�k�9�o�9�l�9n�9n�9�k�9�i�9n�9�m�9Ym�9�n�9�p�9�m�9�l�9n�9x   x   ol�9xj�9�m�9Jm�9�n�9<n�9�n�9-r�9�m�9�m�95r�9�m�9�n�9�q�95n�9�n�9�m�9m�9om�9k�9�l�9ol�9$o�9�i�9�n�94r�9�l�9�j�9p�9hl�9x   x   �m�9�n�9�o�9.i�9en�9Ul�9�l�9�k�9Nj�9(m�9�m�9�i�9qk�9�l�9�l�9�n�9�i�9	q�9�m�9�l�9Nn�9�n�9�n�9+n�9�o�9tp�9o�9nm�9�m�9�n�9x   x   �k�9�n�9�o�9�m�9p�9�p�9�k�9k�9�n�9�k�9�n�9ok�9�k�90p�9�n�9bn�9n�9o�9[m�9fo�9�m�9�j�9�p�9rr�9Qh�9_r�98p�9�l�9�m�9�n�9x   x   yk�9om�9�q�9k�9o�9�p�9Mm�9vq�9`m�9m�9�q�9�l�95p�9Fp�9Tk�9r�9!n�9�j�9�k�9�k�9�n�9�j�9�o�9n�9am�9�o�9$j�9�l�9�l�9pm�9x   x   �n�9�n�9m�9�k�9yo�9}l�9�n�9n�9�n�9zn�97n�9�l�9�n�9Tk�9�k�9o�96n�9�n�9�o�9�o�9&o�9im�9�l�9�l�9�m�9�m�9�o�9Aq�9�m�9�m�9x   x   )n�9o�9�p�9�n�95n�9Pn�9�k�9-o�9�n�9�k�9�n�9�n�9dn�9r�9	o�9xm�9�o�9Im�9�n�9n�9�n�9�n�9�l�9�l�9�m�9|n�9+m�9kn�9;o�9�n�9x   x   �m�9cn�9o�9vi�9�n�9Qo�9�p�9�p�9q�9�o�9�m�9�i�9n�9"n�9:n�9�o�9?r�9�l�9(l�9tm�9hm�9�j�9�k�9�k�9}n�9�m�9�l�9�l�9�q�9�o�9x   x   kk�9�n�98p�9�l�9l�9�m�91m�9Gm�96m�9�l�9m�9q�9o�9�j�9�n�9Im�9�l�9�p�9o�9�m�9n�9Xp�9No�97m�9�l�9To�9Sp�9,l�9�n�9n�9x   x   �l�9�m�9�n�9�m�9@l�9$o�9�p�9^o�9�k�9n�9om�9�m�9]m�9�k�9�o�9�n�9+l�9o�9�k�9�o�9n�9�o�9io�9[p�9=l�9�n�9�m�9�m�9�n�9l�9x   x   �m�9Vj�9cm�9�o�9`n�9|m�9m�9mo�9�o�9�m�9!k�9�l�9jo�9�k�9�o�9n�9qm�9�m�9�o�9n�9�n�9wn�9	m�9�o�9�m�9�l�9}m�9�p�9m�9�n�9x   x   Wl�9l�9�l�9Rl�9zm�9�i�9�l�9�k�9Nl�9�k�9�l�9Qn�9�m�9�n�9*o�9�n�9gm�9n�9n�9�n�9�w�9o�9Do�9�m�9Zn�9Ho�9yo�9m�9Em�9=o�9x   x   �j�9�o�9�j�9�o�9�o�9aq�9p�9:k�9	p�9�i�9ql�9�n�9�j�9�j�9gm�9�n�9�j�9Wp�9�o�9zn�9o�9!o�9�o�9�j�9;n�9�l�9k�9Yl�9�n�9kk�9x   x   �p�9�m�9Yj�9kn�9�k�9�l�9�i�9�l�9'r�9n�9$o�9�n�9�p�9�o�9�l�9�l�9�k�9Ro�9lo�9m�9Go�9�o�9�l�9�l�9,n�9�o�9�o�9�m�9	p�9cn�9x   x   �o�9�m�9m�9�n�9_o�9�n�9�n�9�n�9�n�9�m�9�i�9+n�9qr�9n�9�l�9�l�9�k�9:m�9]p�9�o�9�m�9�j�9�l�9�l�9$m�9�r�9�n�9[j�9m�9Fo�9x   x   �n�9�o�9�p�9fq�94p�9�m�9�o�9�k�9fj�9Xm�9�n�9�o�9Rh�9fm�9�m�9�m�9~n�9�l�9=l�9�m�9Yn�9<n�9/n�9m�9i�9mo�97n�9�l�9�j�9�k�9x   x   �p�96o�9]m�9m�9�p�9'q�9p�9�n�9-q�9�n�97r�9xp�9Zr�9�o�9�m�9yn�9�m�9So�9�n�9�l�9Eo�9�l�9�o�9�r�9no�9�r�9�o�9�q�9n�9q�9x   x   ]o�9m�9ej�9�l�9rn�9n�9Sl�9n�9Zm�9�p�9�l�9o�99p�9"j�9�o�9'm�9�l�9Rp�9�m�9|m�9yo�9k�9�o�9 o�9=n�9�o�9l�9hn�9tl�9�m�9x   x   �o�9Qq�9r�9�o�96k�9�k�9�o�9n�9�o�9�m�9�j�9om�9�l�9�l�9Eq�9ln�9�l�90l�9�m�9�p�9m�9Xl�9�m�9Xj�9�l�9�q�9gn�9�o�9Pk�9�j�9x   x   �l�97k�9l�9�m�9�j�9�j�9�l�9�o�9k�9�l�9p�9�m�9�m�9�l�9�m�9;o�9}q�9�n�9�n�9m�9@m�9�n�9
p�9m�9�j�9
n�9tl�9Rk�9/l�95m�9x   x   �l�9tm�9Pk�9-m�9�l�9�m�9o�9�k�9,o�9n�9nl�9�n�9�n�9qm�9�m�9�n�9�o�9n�9�l�9�n�9@o�9mk�9an�9Eo�9�k�9q�9�m�9�j�94m�9�k�9x   x   ˍ�9	��9>��9m��9K��99��9ی�9֑�9��9Ó�9�9��9͒�9���9���9z��9���9��9H��9���9��9V��9���9`��9���9���9���99��9X��9���9x   x   
��9���9���9ْ�9��9/��9J��9���9���9F��9���9,��9���9Ѝ�9���9���9���9��9��9��9���9���9���9���9Č�9���9.��9���9?��9���9x   x   ?��9���9U��9
��9A��9I��9e��9w��9X��9-��9̓�9���9͑�9���9��9t��9:��9A��9���9'��9/��9"��96��9��9��9��9���9r��9���9,��9x   x   g��9ڒ�9��9���9��9��9���9z��9���9���9���9���9Г�9���9��9��9$��9���9���9���9���9~��9{��9j��9���9Ք�9[��9{��9���9ґ�9x   x   G��9��9>��9��9��9���9���9���9/��9���9���9Y��9���9���9y��91��9���9��9���9_��9x��9ϐ�9p��9��9��9Տ�9��9$��9���9��9x   x   9��9/��9G��9 ��9���94��9���9���9���9���9���9~��9���9���9���9���9@��9Փ�9l��9���9���9���9��9���9��9U��9���9���9{��9;��9x   x   ،�9L��9b��9���9���9���9��9���9Ȍ�9>��9w��9���9��9��9e��9��92��9o��9i��9:��9���9T��9S��9ϔ�9 ��9a��9 ��9���9U��9P��9x   x   ۑ�9���9w��9|��9���9���9���9*��9l��9���9���9.��9��9��9'��9��9���9��9���9ɏ�9���9���9���9Œ�9���9;��9���9$��9���9b��9x   x   ��9���9U��9���92��9���9ǌ�9l��9���9Ƒ�9h��9n��9��9��9���9��9Q��9��9e��9W��9���9Đ�9���9���9���9r��9��9���9 ��9R��9x   x   ē�9C��9)��9���9���9���9;��9���9ɑ�9��91��9ʐ�9Ƒ�9��9���9���9R��9��9��9ߑ�9��9
��9%��95��9���9]��9J��9���9���9$��9x   x   ĕ�9���9̓�9���9���9���9u��9���9i��91��9(��9A��9���9��9��9Θ�9���9V��9<��9m��9���9���9Y��9���9 ��9��9.��9���9n��9��9x   x   ��9-��9���9���9[��9���9���9+��9k��9̐�9D��9>��9%��9��9f��9U��9��9���9��9ǐ�9 ��9��9��9G��9v��9%��9���9ҏ�9���9���9x   x   Β�9���9͑�9͓�9���9���9ߓ�9ߒ�9��9�9���9%��9���9��9*��9���9B��9a��9���9���9��9���9��9���9ӓ�9M��9���9���9��9���9x   x   ���9̍�9���9���9���9���9��9��9��9��9��9��9��9���9��9C��9���9V��9Ƒ�9U��9X��9̓�9���9ђ�9���9T��9
��95��9���9ʒ�9x   x   ���9��9��9��9w��9���9`��9(��9���9���9��9c��9+��9��9��9��9��9Ґ�9���9G��9_��9���9���92��9c��9;��9���9��9s��9^��9x   x   |��9���9x��9��91��9���9���9��9���9���9̘�9S��9���9E��9��9v��9���9T��9���9L��9���9*��9��99��9t��9���9��9x��9���9���9x   x   ���9���9:��9"��9���9C��93��9���9T��9V��9���9��9B��9���9ߑ�9���9G��9q��9��9R��9���9.��9���9b��9$��9=��9W��9&��9��94��9x   x   
��9��9@��9���9��9ӓ�9n��9��9��9��9U��9���9]��9T��9͐�9V��9p��9��9D��9֓�9��9{��9ܐ�9���9;��9e��9��9���9���9?��9x   x   I��9��9���9���9���9m��9l��9���9d��9��9@��9��9���9ɑ�9���9���9��9C��9���98��9Ց�9���9���9���9 ��9���9��9ד�97��9��9x   x   ���9��9 ��9���9d��9���98��9ʏ�9T��9ݑ�9j��9Đ�9���9W��9C��9K��9U��9ד�98��9C��9��9
��9q��9��9��9��9J��9y��9F��9��9x   x   ��9���9+��9���9v��9���9���9���9���9��9���9 ��9��9X��9\��9���9���9��9Ց�9��9u��9��9���9v��9ڒ�9���9(��9���9ڑ�9���9x   x   Y��9��9$��9���9ϐ�9���9W��9���9̐�9��9���9��9���9͓�9���9*��9+��9~��9���9��9��9m��9��9���9��9"��9���9���9֏�9��9x   x   ���9���9/��9x��9n��9��9O��9���9���9&��9U��9��9��9���9���9��9���9ې�9~��9n��9��9��9֓�9��9��9���9.��9h��9ԑ�9��9x   x   f��9���9��9k��9��9���9ϔ�9ƒ�9���93��9���9D��9���9Β�9-��9>��9^��9���9���9��9s��9���9��9��9��90��9*��9%��9��9B��9x   x   ���9Ȍ�9��9���9#��9��9 ��9���9���9���9��9v��9ѓ�9���9`��9q��9$��99��9��9��9ג�9��9��9��9���9��9ޏ�9W��9���9���9x   x   {��9���9��9Д�9ӏ�9R��9a��99��9r��9Z��9��9$��9J��9X��9@��9���9@��9d��9Ð�9��9���9%��9���93��9��9���9��9t��9���9���9x   x   ���92��9���9^��9��9���9#��9���9��9D��9+��9���9���9	��9���9��9X��9��9��9G��9+��9���9-��9(��9؏�9��9���9;��9r��9��9x   x   5��9���9n��9}��9$��9���9���9&��9���9���9���9֏�9���96��9���9w��9)��9��9ד�9x��9���9���9g��9#��9V��9t��9:��9���9P��9=��9x   x   Y��9C��9���9���9���9x��9W��9���9 ��9���9m��9���9
��9���9u��9���9��9���9:��9C��9ܑ�9׏�9ԑ�9��9���9���9s��9S��9ʔ�98��9x   x   ��9���9)��9Б�9~��9:��9S��9b��9T��9$��9
��9���9���9͒�9]��9č�98��9D��9��9��9���9���9��9B��9��9���9��9<��94��9���9x   x   z��9���9׶�9���9}��9���9۹�9C��9��9s��9���9ٸ�9��9��9¸�9���9���9��9��9��9���9��9Ѹ�9��9��9޺�9���9M��9���9g��9x   x   ���9��96��9��9���9U��9	��9��9Ҵ�9t��9���9ֵ�9���9{��9���9���9���9B��9}��9���9(��9��9���9{��9O��9���9���9r��9��9���9x   x   ׶�99��9��9&��9���9��9ٳ�9���9O��9[��9o��9[��9��9��9T��9:��99��9��9q��9ϵ�9G��9E��9ɴ�9Ų�91��9]��9���9v��9+��9��9x   x   ���9��9 ��9`��9��9��9z��99��9���9���9*��9���9��9c��9��9y��9Ӻ�9[��9۴�9ȶ�9��9��9��9��9��9��9��96��9o��9Դ�9x   x   ���9���9���9!��93��9���9���9���9���9���9��9G��9��9ַ�9߹�9���9���9��95��9��9õ�9I��9Ÿ�9��9q��9��9ܳ�9���9<��9���9x   x   ���9T��9���9��9���9���9e��9%��9@��9��9��9���9.��9f��9���9C��9��9���9��9���9��9´�9���9_��9��9���95��9Դ�9��9f��9x   x   ܹ�9��9ٳ�9{��9���9b��9׸�9���9]��9���9R��9O��9d��9_��9$��9���9!��9K��9X��9��9E��9��9��9���9��9��9���9ں�9ٷ�9���9x   x   @��9��9���95��9���9%��9���93��9	��9��9���9��9���9ò�9��9���9P��9���95��9��9���9���9b��9���9��9\��9E��9ܸ�9j��9���9x   x   ��9Դ�9S��9���9���9?��9_��9��9A��9d��9��9��9��9���9ĸ�9k��9G��9���9 ��9��9N��9w��9���9ȷ�9k��9,��9��9&��9��9h��9x   x   r��9w��9^��9���9���9��9���9��9j��9յ�9���9��97��9���9��9���9��9���9w��9
��9ǳ�9���9u��9���9a��9+��9��9��91��9ַ�9x   x   ���9���9o��9)��9{��9���9U��9���9��9���9@��9���9v��9&��9۲�9���9���9G��9Գ�9#��9ΰ�9���9���9���9���9��9��9��9i��9���9x   x   Ӹ�9ֵ�9Y��9���9D��9���9U��9��9��9 ��9���9���9���9��9���9u��9���9��9Ŷ�9*��9ȴ�9��9Ҷ�9k��9���99��9k��9}��9_��9&��9x   x   ��9���9��9	��9��9-��9k��9���9"��9;��9x��9���9��9]��9	��9���9���9���9J��9.��9���9~��9���9��9���9��9���9>��9 ��9&��9x   x   ��9{��9��9f��9ҷ�9c��9a��9���9���9~��9&��9��9X��9��9T��9��9��9ø�9��9ҷ�9ǳ�9;��9I��9��9ҷ�9p��9ٷ�9_��9��9��9x   x   ���9���9S��9��9۹�9���9'��9��9���9��9۲�9ö�9��9R��9���9Q��9Զ�9���9���9��9`��9���9��9��9���9w��9���9��9ڶ�9���9x   x   ���9���99��9y��9���9B��9���9���9k��9���9���9x��9���9��9S��9p��9i��9[��9���9&��9���9`��9���9۳�9-��9���9��9���9[��9���9x   x   ���9���98��9ֺ�9���9��9!��9L��9E��9��9���9���9���9��9׶�9i��9���9g��9h��9n��92��9���9���9K��9���9��9��9)��9��9C��9x   x   ��9B��9��9X��9���9���9N��9���9���9���9D��9��9���9Ǹ�9Ŷ�9[��9g��9��9E��9G��9q��9���9ɵ�9���9ϵ�9'��9ĸ�9n��9O��9���9x   x   ��9��9q��9ܴ�94��9��9W��94��9���9{��9ҳ�9ȶ�9I��9��9���9���9f��9E��9J��90��9���9��9}��9V��9��9��9���9Ƶ�9���9���9x   x   ��9���9ҵ�9ʶ�9��9���9��9��9��9��9#��9/��9'��9շ�9��9'��9n��9H��91��9j��9��9t��9��9���9c��9���9ȸ�9ƴ�9��9K��9x   x   ���9,��9H��9��9ŵ�9!��9J��9���9L��9ĳ�9Ӱ�9˴�9���9ʳ�9a��9���91��9l��9���9��9/��9��9��9��9ٳ�9]��9T��9޲�9|��9��9x   x   ��9��9D��9��9H��9´�9��9���9u��9���9���9���9{��99��9���9^��9���9ô�9��9t��9��9���9���9���9,��9���9Ƿ�9m��9���9д�9x   x   ͸�9���9ʹ�9#��9Ÿ�9���9#��9e��9���9u��9���9̶�9���9J��9~��9���9���9ɵ�9���9��9���9���9���9���9���9���9q��9���9ʳ�9���9x   x   ��9{��9Ų�9��9��9\��9���9���9ŷ�9���9���9j��9!��9��9#��9߳�9O��9���9U��9���9��9���9���9ش�9��9b��9���9+��9/��9ض�9x   x   ��9M��9.��9��9o��9��9��9��9k��9`��9���9���9���9շ�9���9*��9���9е�9��9a��9ݳ�9*��9���9"��9��9��9���9A��93��9��9x   x   ��9���9[��9���9��9���9��9\��9+��9.��9��97��9��9q��9w��9���9��9)��9��9���9]��9���9���9c��9��9���9���9+��9���9ٶ�9x   x   ���9���9���9��9س�97��9���9D��9��9��9 ��9n��9���9Է�9���9��9��9���9���9Ǹ�9R��9Ʒ�9m��9���9���9���9��9ٸ�9��9O��9x   x   J��9s��9r��96��9���9ִ�9غ�9ڸ�9'��9��9��9y��9@��9a��9��9���9*��9l��9ʵ�9ƴ�9ݲ�9n��9���92��9A��9.��9ٸ�9��9���9H��9x   x   ���9��9(��9m��9<��9��9ط�9k��9��91��9k��9[��9��9��9ض�9V��9��9J��9���9��9��9��9ɳ�9+��92��9���9��9���9���9(��9x   x   c��9���9��9Ѵ�9���9h��9���9ö�9g��9ѷ�9���9(��9#��9��9���9���9D��9���9���9Q��9��9Ѵ�9���9׶�9��9ض�9P��9F��9(��9Ӹ�9x   x    ��9J��9���9���9���9_��9���9��9���9D��9���9T��9���9:��9���9���9���9���9$��9o��9n��9���9���9���9���9z��9��9f��9��9��9x   x   Q��9f��9���9a��9���9N��9���9���9���9��9���9j��9���9���9W��9���9@��9���9	��9P��9��9?��9���93��97��9r��9!��9y��9��9M��9x   x   ���9~��9\��9���9��9���9=��9���9R��9��9���9|��9���9���9���9t��9���9���9`��9���9���9���9��9���92��9f��9j��9\��93��9W��9x   x   ���9_��9���9���9���9(��9���9&��9��9s��95��9���9���9���9l��9���9��9V��9���9Q��9���9���9���9���9���9O��9���9_��9���9���9x   x   ���9���9��9���9/��9���9s��9^��9��9q��9���9��9G��9���9��9q��9���9
��9���9x��9y��9���9��9���9P��9���9<��9��9��9z��9x   x   Z��9K��9���9%��9���9���9F��9���9��9p��9���9���9���9X��91��9��9���9u��9���9K��9���9
��9'��9`��9���9~��9��9���9Y��9���9x   x   ���9���9<��9���9u��9G��9���9��9���9���9���9��9���9���9S��9��9S��9���9$��9���9b��9���9���96��9���9���9���9g��9��9D��9x   x   ��9���9���9#��9_��9���9��9���9���92��9��9_��9��9j��9���9s��9���9���9A��9��9��9���9��9���9���9)��9��9Z��9K��9���9x   x   ���9���9U��9��9
��9��9���9���9"��9%��9c��9���9M��9���9���9T��9��9v��9���9���9���9	��9���9���9p��9>��9z��9���9���9���9x   x   D��9���9��9t��9r��9s��9���90��9"��9R��9���9���9m��9:��9���9��9m��9y��9���9���99��9?��9q��9���9���9���9��9��9/��9���9x   x   ���9���9���94��9���9���9���9��9b��9���9P��9���9��9|��9���9_��9���9v��9���9���9���9���9A��9���9���9���9���9<��9|��9P��9x   x   U��9n��9|��9���9��9���9��9[��9���9���9���9���9���9F��9���9L��9���9���9N��9I��9���9��9e��9���90��9��9���9��9��9���9x   x   ���9���9���9���9K��9���9���9��9J��9q��9��9���9��9��9}��9V��9���9���9��9:��9 ��9���9b��9(��9��9���9l��9���9a��9���9x   x   =��9���9���9���9���9W��9���9d��9���9>��9{��9G��9��9��9v��9>��9z��9m��9���9���9c��9A��9��97��9��9*��9���92��9i��9���9x   x   ���9\��9���9k��9��91��9U��9���9���9���9���9���9���9x��9]��9��9���9���9X��9j��9���9u��9���9���9 ��9���9���9���9?��99��9x   x   ���9���9s��9���9r��9��9	��9s��9Y��9��9Y��9I��9Y��9@��9��9���9���9���9��9`��9���9���9��9���9���98��9��9{��9���9.��9x   x   ���9A��9���9��9���9���9R��9���9��9h��9���9���9���9u��9���9���9���9-��9���9���9Z��9F��9	��9���9��9���98��9���9Y��9*��9x   x   ���9���9���9V��9��9t��9���9���9w��9{��9v��9���9���9i��9���9���9-��9a��9c��9���9h��9���9���9Q��9��9���9��9.��9���9b��9x   x   "��9
��9[��9���9���9���9$��9@��9���9���9���9M��9��9���9W��9��9���9e��9���9��9"��9>��9���9-��92��9/��94��9��9>��9���9x   x   o��9N��9���9Q��9w��9Q��9���9~��9���9���9���9G��9:��9���9i��9`��9���9���9"��9q��9+��98��9���9,��9p��9���9 ��9N��9%��9&��9x   x   n��9��9���9���9x��9���9c��9��9���9;��9���9���9��9b��9���9���9[��9d��9#��9-��9e��9��9���9��9.��9��9p��9M��9:��9p��9x   x   ���9;��9���9���9���9��9���9���9��9B��9���9��9���9?��9x��9���9O��9���9<��97��9��9v��9#��9b��9d��9%��91��9I��9<��9��9x   x   ���9���9��9���9��9+��9���9!��9���9u��9D��9f��9a��9��9���9��9��9���9���9���9���9#��9���9��9g��9	��9���9���9���9��9x   x   ���93��9���9���9���9b��95��9���9���9���9���9���9%��94��9���9���9���9N��9,��9*��9��9\��9��9{��9��9���9���9���9���9���9x   x   ��95��93��9���9M��9���9���9���9o��9���9���92��9��9��9��9���9��9��90��9q��9.��9b��9h��9��9���9]��9/��9���9���9k��9x   x   y��9p��9h��9Q��9���9���9���9,��9?��9���9���9��9���9'��9���96��9���9���9/��9���9��9&��9	��9���9^��9���9���9O��9���9���9x   x   ��9!��9g��9���97��9��9���9��9x��9��9���9���9n��9���9���9��96��9��94��9��9q��96��9���9���9/��9���9���9h��9_��94��9x   x   k��9z��9^��9f��9��9���9h��9Z��9���9��99��9��9���9/��9���9|��9���9-��9
��9N��9J��9J��9���9}��9���9M��9f��9R��9���9���9x   x   ��9~��92��9���9 ��9X��9��9P��9���9/��9���9��9_��9k��9?��9���9[��9���9>��9#��95��9<��9���9���9���9���9]��9���9/��9���9x   x   ��9H��9W��9���9y��9���9B��9���9���9���9T��9���9���9���9?��9+��9*��9f��9���9'��9o��9��9��9���9k��9���98��9���9���9���9x   x   ���9��9m�9���9�9��9��9��9��9��9	�9��9h�9��9��9	�9��9?�9��9��9O	�9��9���9w�9N�9��9�9' �9(�9Q�9x   x   ��9H�9@�9��9@�9��9/�9��91�9a�9) �9��9��9o�9Y�9��9q�9��9��9���9��9��9� �9�9��9��9"�9��9�	�9 �9x   x   n�9>�96�9#�9��9J	�9k�9_�9�9  �9��9,�9��9��9� �9;�9��9�9��9���9�9�9��9��9��9��9�99�9�9��9x   x   ���9��9&�9� �9�9��9� �9��9� �9�9��9��9b�9��9�9 	�9��9��9��9��92�9���9?�9��9���9&�9��9���9��97�9x   x   �9A�9��9�9l�9��9��9��9��9��9?�9%�9��9{�9X�9O�9e�9��9�9�9n�9	�9a�9��9��9.�9�9���9��9o��9x   x   ��9��9H	�9��9��9-�9��9��94�9��9x�9; �9��9��9� �9��9I�9��9v�9��9 �9r�9�97	�9��9a�9��9m�9!�9�9x   x   ��91�9k�9� �9��9��9c�9��9��9��9��9���9A�9���9D�91�9D�9��9)�9��9��9� �92�9�9��9��9��9��9��9�9x   x   ��9��9\�9��9��9��9��9��90�9��9��9U�95�9��9%�9��9��9��9��9��9Y�9��9?�9?�9��9��97�9B�9��9"�9x   x   ��93�9�9� �9��95�9��93�93�9��9D�9��9"�9;�9��9��9l�9�9��9� �9�9� �9���9��93�9~�9�9��9�9�9x   x   ��9]�9���9�9��9��9��9��9��9��9� �9��9��9��95�9�9� �9��9��9��9��9��9��9�9�9��9��9�9��9*�9x   x   	�9% �9��9��9=�9y�9��9��9D�9� �9���9�9�9.�9��9�	�9��9��97�9" �9��9��9��9��9<�9��9w�9��9��9��9x   x   ��9��91�9��9%�9> �9���9V�9��9��9�9��9��9[ �9���9��9��9;�9��9�9�9v �9>�9|�9��9;�9s�9=�9� �9��9x   x   f�9�9��9c�9��9��9A�99�9!�9��9�9��9��9C�9&�9@�9��9 �9%�9>�9��9��95�9��9��9��9��9��9��9��9x   x   ��9k�9��9��9y�9��9���9��9:�9��9.�9] �9C�9��9��9��9��9h�9��9�9K�9��9��90�9.�9��9��9��9b�9��9x   x   ��9X�9� �9�9U�9� �9A�9"�9��91�9��9���9$�9��9$�9W�9��9�9��9O�9��9��9�9�9T�90�9��9Z�9  �9��9x   x   
	�9��9@�9	�9O�9��91�9��9��9�9�	�9��9B�9��9W�9��9��9��98�9
�9��9M�9��9Y�9��9�9��9r�9X�96�9x   x   ��9q�9��9��9f�9J�9G�9��9m�9� �9��9��9��9��9��9��9� �9��9��9��9��9��9��9�9��94�9�9G�9��9��9x   x   @�9��9�9��9��9��9��9��9	�9��9��98�9�9j�9�9��9��9+�9$�9��9E�9R�97�9��9��9�9�9H�9��9�9x   x   ��9��9��9��9�9y�9&�9��9��9��9;�9��9)�9��9���98�9��9#�9��9��9-�94�9��9��9��9�9��9 �9c �9g�9x   x   ��9���9���9��9�9��9��9��9� �9��9% �9�9C�9�9N�9	�9��9��9��9&�9]�9+�9��9��9�9��9;�94�9��9u�9x   x   Q	�9��9�95�9l�9�9��9Z�9�9��9��9�9��9G�9��9��9��9A�9-�9]�9��9B�9��9�9�9��9��9F�9�9E�9x   x   ��9��9�9���9�9w�9� �9��9� �9��9��9t �9��9��9��9J�9��9Q�92�9+�9D�97�9��9�9�9O�9	�9��9���9��9x   x   ���9� �9��9>�9e�9�9,�9<�9���9�9��9?�98�9��9�9��9��99�9��9��9��9��9��9��9��9��9v�9�9��9�9x   x   w�9�9��9��9��9:	�9�9B�9��9�9��9x�9��92�9�9[�9�9��9��9��9�9�9��9��9��9{�9�9��9��9�9x   x   N�9��9��9���9��9��9��9��92�9�9=�9��9��90�9S�9��9��9��9��9�9�9�9��9��9��9l�9&�9��9x�94�9x   x   ��9��9��9"�9,�9`�9��9��9��9��9��9;�9��9��9.�9�97�9�9��9��9��9N�9��9}�9m�9��9m�9/�9�9��9x   x   �9%�9�9��9�9��9��95�9�9��9w�9s�9��9��9��9��9�9�9��9<�9��9�9v�9�9%�9m�9�9D�9��9 �9x   x   & �9��97�9���9���9l�9��9B�9��9�9��9?�9��9��9X�9p�9E�9F�9��95�9K�9��9�9��9��9/�9F�9��9�9���9x   x   '�9�	�9�9��9��9�9��9��9�9��9��9� �9��9d�9" �9[�9��9��9a �9��9!�9���9��9�9x�9�9��9�9#�9��9x   x   X�9 �9��98�9r��9�9�9 �9�9+�9��9��9��9��9��92�9��9�9d�9p�9F�9��9�9�90�9��9��9���9��9,�9x   x   4�9e-�9"/�9j/�9
.�9�-�9.*�9P+�9�2�9.�9L+�9�,�9;)�9�*�9�,�9*�9h,�9H)�9)�9i,�9`,�9.�9�2�9�+�9
+�9N.�9�-�9I/�9�-�9O-�9x   x   c-�96*�95,�9b)�9�-�9e0�9�)�9�.�9-�9�+�9f0�9�.�9a.�96-�9s-�9�-�9Z.�9G/�9�.�9�/�9E+�9h-�9�-�9�*�9/�9�,�9E*�9�,�9y+�9�,�9x   x   !/�94,�9�-�9+�9�)�9G*�9B+�9�.�9�+�9p0�9�,�9�,�9-�9+�9?-�9*�9,�9Z,�9�-�9�0�9�+�9�/�9"+�9�)�9�+�9�+�9,�9�+�9�.�9�+�9x   x   l/�9a)�9+�9�+�9/�9W+�95.�9�.�9�-�9/�9�-�9�/�9:-�9$+�9A,�95.�9]0�9W-�9�-�9!.�9�-�9M.�9�+�9�.�9�)�9�+�9/+�9�.�9d.�9�-�9x   x   .�9�-�9�)�9/�9G2�9",�9�-�9�*�9�+�9�-�92-�9|+�9�+�9�)�9}*�9�*�9-�9_.�9*,�9s+�99.�9�+�9�2�9Y/�9s+�9�,�9e-�9�/�9�0�9/�9x   x   �-�9g0�9I*�9\+�9,�9+,�9�-�9�,�9/�9G,�9�,�9�.�9#/�9w/�9�/�9�,�9�+�9D/�9�+�9Z-�9f,�9�+�9#+�9 *�9x/�9�.�9�*�9�*�9e,�99*�9x   x   **�9�)�9?+�92.�9�-�9�-�9-�9�,�9�.�9�.�9k2�9�,�9�)�9�,�9}1�9�/�9Y.�9�,�9.�9}-�9).�9u.�9x+�9�)�9~+�9�+�9G,�9X.�9+�9&-�9x   x   O+�9�.�9�.�9�.�9�*�9�,�9�,�9�)�96+�9I,�9�+�9�,�99,�97,�9,�9+�9*�9�+�9�,�9�*�9�.�9x.�92/�9	+�9�,�9�)�9�,�9�,�9�)�9Z-�9x   x   �2�9-�9�+�9�-�9�+�9/�9�.�97+�9&,�9,�9-�9�-�9?-�9�,�9�+�9e+�9�.�9/�9�,�9�-�9,�9-�9m2�9�-�9�-�9<,�9�,�9s-�9�+�9B.�9x   x   .�9�+�9u0�9/�9�-�9E,�9�.�9F,�9 ,�9�/�9�/�9_0�91.�9�+�9�,�9*.�9�,�92-�9�.�9�/�9�+�9�-�9�0�9#)�9<*�9m.�9z,�9;+�9�*�9�/�9x   x   J+�9j0�9�,�9�-�93-�9�,�9f2�9�+�9-�9~/�9�3�9�/�9�.�9�+�9m2�9�,�9H-�9�-�9�-�9�0�9�+�9,�9.�9�,�9B,�9=/�9�,�9k+�9S-�9�,�9x   x   �,�9�.�9�,�9�/�9z+�9�.�9~,�9�,�9�-�9a0�9�/�9|-�9�+�9d,�9v/�9�*�9�/�9p,�9p.�9E,�9a/�9�.�9�-�9E.�90*�9�*�9�-�9�.�9�/�9U.�9x   x   >)�9d.�9-�9<-�9�+�9'/�9�)�97,�9A-�94.�9�.�9�+�9�+�9�.�9�+�9G-�9(-�9�.�98*�9 .�9�/�9�.�9�-�9^-�9t*�9�,�9D.�9&-�9�/�9�.�9x   x   �*�94-�9+�9'+�9�)�9z/�9},�95,�9�,�9�+�9�+�9c,�9�.�9�)�9d+�9�*�9F-�9�)�9(+�9�/�9]'�9E,�9�-�9p.�9�.�9�-�9V,�9�(�99/�9�*�9x   x   �,�9t-�9:-�9A,�9|*�9�/�9z1�9,�9�+�9�,�9m2�9w/�9�+�9a+�9a-�9�-�9�-�9+�9�-�90�9Q-�9d0�9,�9�,�9<,�9�/�90-�9�.�9 .�9i+�9x   x   *�9�-�9 *�98.�9�*�9�,�9�/�9"+�9e+�9+.�9�,�9�*�9L-�9�*�9�-�9)�9-�9�.�9*-�9O/�9o.�9--�9-�9�,�9�-�9�.�9�/�9M.�9�-�9�,�9x   x   j,�9V.�9,�9_0�9-�9�+�9Y.�9*�9�.�9�,�9F-�9�/�9(-�9D-�9�-�9-�9�/�9(-�9�+�9�,�9�,�9�0�9�0�9c0�9T,�9d,�9�*�9�,�9�0�9�,�9x   x   H)�9H/�9[,�9U-�9\.�9E/�9�,�9�+�9/�9.-�9�-�9s,�9�.�9�)�9+�9�.�9)-�9J,�9".�9<.�9�/�9c,�97-�9�/�9�.�9�.�9�,�9 -�9�-�9,�9x   x   )�9�.�9�-�9�-�9-,�9�+�9.�9�,�9�,�9�.�9�-�9p.�93*�9&+�9�-�9(-�9�+�9!.�9�+�9-�9�,�9�-�9�+�9�,�9?+�9�-�9+�9�-�9�-�9!+�9x   x   g,�9�/�9�0�9$.�9s+�9[-�9�-�9�*�9�-�9�/�9�0�9E,�9�-�9�/�90�9N/�9�,�9<.�9
-�9+�98.�9H.�9�+�9�-�9s.�9
-�9f/�9�/�9.�9�/�9x   x   _,�9F+�9�+�9�-�9<.�9i,�9+.�9�.�9,�9�+�9�+�9b/�9�/�9b'�9S-�9o.�9�,�9�/�9�,�97.�9|+�9.�9c+�9�/�9",�9.�9�,�98)�9�/�9;.�9x   x   .�9i-�9�/�9L.�9�+�9�+�9z.�9w.�9-�9�-�9,�9�.�9�.�9@,�9_0�9.-�9�0�9d,�9�-�9I.�9#.�9s.�9-�91�9[-�91�9c+�9�-�92/�9Y,�9x   x   �2�9�-�9$+�9�+�9w2�9+�9{+�93/�9k2�9�0�9.�9�-�9�-�9�-�9,�9-�9�0�99-�9�+�9�+�9a+�9-�9�/�9(-�9+�9n.�9.�9�.�9?.�9�/�9x   x   �+�9�*�9�)�9�.�9X/�9�)�9�)�9+�9�-�9()�9�,�9E.�9b-�9k.�9�,�9�,�9`0�9�/�9�,�9�-�9�/�91�9%-�9�-�9�.�9�,�9�-�9�*�9`*�9~.�9x   x   	+�9/�9�+�9�)�9r+�9t/�9+�9�,�9�-�9;*�9C,�9/*�9s*�9�.�9<,�9�-�9V,�9�.�9;+�9v.�9",�9[-�9+�9�.�9L*�9+�9�-�9�*�9�,�9�+�9x   x   N.�9�,�9�+�9�+�9�,�9�.�9�+�9�)�9<,�9l.�9?/�9�*�9�,�9�-�9�/�9�.�9b,�9�.�9�-�9-�9}.�91�9r.�9�,�9+�92-�9�-�9�+�9r+�9�,�9x   x   �-�9C*�9",�9.+�9g-�9�*�9I,�9�,�9�,�9y,�9�,�9�-�9@.�9S,�92-�9�/�9�*�9�,�9!+�9i/�9�,�9e+�9.�9�-�9�-�9�-�9�-�9t,�9*�9+�9x   x   G/�9�,�9�+�9�.�9�/�9�*�9Z.�9�,�9s-�98+�9l+�9�.�9#-�9�(�9�.�9P.�9�,�9-�9�-�9�/�97)�9�-�9�.�9�*�9�*�9�+�9v,�9q/�9�+�9/�9x   x   �-�9x+�9�.�9c.�9�0�9f,�9+�9�)�9�+�9�*�9S-�9�/�9�/�9:/�9�-�9�-�9�0�9�-�9�-�9.�9�/�91/�9;.�9Y*�9�,�9p+�9*�9�+�9�/�9}.�9x   x   K-�9�,�9�+�9}-�9/�96*�9(-�9X-�9>.�9�/�9�,�9Y.�9�.�9�*�9j+�9�,�9�,�9,�9'+�9�/�9<.�9Y,�9�/�9y.�9�+�9�,�9�*�9/�9y.�9.,�9x   x   rX�9�V�9�T�9X�9JW�9T�9�W�9tV�9�T�9�V�9.T�9�W�9�W�9�W�9�V�9�T�9LW�9RV�9�W�9�W�9DU�99W�9�T�9\V�9WW�9�T�9�V�9^W�9�U�9�V�9x   x   �V�9HR�9BY�9�U�9qT�9aX�9�Z�9�W�9DX�9�X�9-X�9�W�9iZ�9[�9�X�9�X�9[�9#[�9�W�9�W�9QW�9:X�9BW�9�[�9X�9�S�9�V�9�X�9YR�9W�9x   x   �T�9AY�9>Z�9�W�9�X�9iV�9�Z�9�S�9YT�9�W�9�S�9U�9�W�9�U�9x\�9XU�9�W�9,T�9zS�9�X�9WU�9�S�9�Y�9&V�9�Y�9^W�9Z�9{Y�9�T�9 W�9x   x   X�9�U�9�W�9_�9�S�9>X�9rY�9
T�9�Y�9�V�9AV�9�W�9�U�9�Y�9�Z�9�U�9X�9W�9�U�9�Y�9S�99Z�9gX�9S�9�^�9W�9�V�9�W�9�R�9�R�9x   x   JW�9qT�9�X�9�S�9FR�9~X�9PU�9_Y�98V�9�W�9Z�9�V�9�[�9�U�9�Z�9�V�9�Y�9�W�9�V�9�Y�9ZU�9�W�9S�9gS�9�Y�9T�9IV�9�X�9W�9�W�9x   x   T�9aX�9eV�99X�9�X�9�V�9nX�9jV�9�S�9�X�9WR�9oX�91V�9V�9Y�9�R�9XX�9�S�9�U�9�X�9�V�9�W�9HX�9�U�9�W�99U�9�W�9�U�9�W�9�W�9x   x   �W�9�Z�9�Z�9tY�9PU�9mX�9�W�90X�9FZ�9�V�9U�91Y�9V�9IY�9�S�9�W�9RZ�9�X�9,X�9�W�9�V�9sY�9)[�9&[�9�W�9�W�93[�9�T�9�Y�9�X�9x   x   wV�9�W�9�S�9
T�9^Y�9iV�9-X�9bW�9iV�9VW�9Y�9�X�9�X�9�Y�9$W�9�U�93W�9X�9�V�9�X�9GS�9HS�9W�9�V�9�V�9�X�9�V�9�V�9uY�9�V�9x   x   �T�9BX�9UT�9�Y�97V�9�S�9DZ�9eV�9�X�9�X�9W�9`U�9jV�9
Y�9Y�9�V�9:Z�9�R�9�V�9�Y�9rU�9�X�9wT�9T�9]�9~Y�9�U�98Z�9�[�9uT�9x   x   �V�9�X�9�W�9�V�9�W�9�X�9�V�9[W�9�X�9�U�9eT�9iU�9+U�9@X�9KW�9xV�9�Y�9�V�9V�9�W�9�W�9�V�9�S�9hW�9�Y�9�W�9dV�9�Y�9�X�9XS�9x   x   /T�9,X�9�S�9FV�9Z�9VR�9U�9Y�9W�9hT�9�T�9sT�9�W�9'Y�9oU�9rQ�9�Y�93W�9�S�9cX�9U�9&W�9�X�9=Y�9�T�9W�9�U�9�X�9�W�9�W�9x   x   �W�9�W�9 U�9�W�9�V�9qX�91Y�9�X�9aU�9fU�9mT�9!U�9�X�9�X�9<Y�9W�9�W�9�S�9dW�9�W�9�X�9}V�9�T�9�W�9�Y�9�X�9W�9�U�9DW�9tX�9x   x   �W�9jZ�9�W�9�U�9�[�91V�9V�9�X�9iV�9-U�9�W�9�X�9`W�9�U�9�Z�9�U�9�X�9`[�9X�9eV�9GV�9�W�9�W�9�Y�9�W�9�Z�97X�9wV�9U�9JW�9x   x   �W�9[�9�U�9�Y�9�U�9V�9HY�9�Y�9Y�9<X�9(Y�9�X�9�U�9�V�9�Y�9�U�9oZ�9�V�9Y�9�W�9�V�9W�93X�9�U�9HU�9hW�9W�9�X�9�W�9�W�9x   x   �V�9�X�9y\�9�Z�9�Z�9Y�9�S�9&W�9Y�9HW�9qU�9<Y�9�Z�9�Y�9�\�9�X�9�W�9[�9)Y�97Y�9X�9�T�9@W�9�Z�9sW�9�U�9�V�9�W�9Z�9[�9x   x   �T�9�X�9WU�9�U�9�V�9�R�9�W�9�U�9�V�9xV�9pQ�9W�9�U�9�U�9�X�9BT�9�Y�9#W�9�R�9�V�9�X�9�W�9�W�9ZX�9lW�9�X�9�W�9S�9�V�9Z�9x   x   GW�9�[�9�W�9X�9�Y�9XX�9QZ�90W�9;Z�9�Y�9�Y�9�W�9�X�9mZ�9�W�9�Y�9EU�9�W�9WX�9�V�9>V�9*X�9NS�9�W�9dV�9�V�9�W�9BW�9HU�9`Y�9x   x   QV�9&[�9(T�9%W�9�W�9�S�9�X�9	X�9�R�9�V�96W�9�S�9b[�9�V�9[�9"W�9�W�9�[�9�W�90X�9�W�9V�92V�9�X�9�W�9�W�9�\�9PX�9�V�9�[�9x   x   �W�9�W�9wS�9�U�9�V�9|U�9.X�9�V�9�V�9V�9�S�9dW�9X�9Y�9)Y�9�R�9YX�9�W�9�W�9�X�9 W�9&Z�9�V�9>X�9�X�9�W�9�V�9PS�9IY�9-Y�9x   x   �W�9�W�9�X�9�Y�9�Y�9�X�9�W�9�X�9�Y�9�W�9gX�9�W�9gV�9�W�92Y�9�V�9�V�91X�9�X�9�V�9�X�9�X�9W�9�X�9iW�9�W�9�W�9�X�9�V�9W�9x   x   EU�9PW�9VU�9S�9\U�9�V�9�V�9FS�9vU�9�W�9U�9�X�9KV�9�V�9X�9�X�9;V�9�W�9�V�9�X�9�S�9�X�9�V�9@X�9 V�9�W�9W�9�X�9eV�9xW�9x   x   =W�9?X�9�S�97Z�9�W�9�W�9sY�9DS�9�X�9�V�9"W�9zV�9�W�9W�9�T�9�W�9)X�9V�9#Z�9�X�9�X�91Z�9RV�9qX�9�W�9jV�9�V�9�U�9IW�9�W�9x   x   �T�9AW�9�Y�9hX�9!S�9MX�9*[�9W�9{T�9�S�9�X�9�T�9�W�96X�9?W�9�W�9NS�91V�9V�9�W�9�V�9QV�9dR�9vX�9�V�9�W�9�X�9�U�91X�9�R�9x   x   ^V�9�[�9"V�9S�9lS�9�U�9%[�9�V�9T�9eW�9<Y�9�W�9�Y�9�U�9�Z�9YX�9�W�9�X�9=X�9�X�9>X�9oX�9uX�9[�9�U�9�Y�9TW�97X�9Y�9�T�9x   x   ]W�9X�9�Y�9�^�9�Y�9�W�9�W�9�V�9]�9�Y�9�T�9�Y�9�W�9JU�9tW�9nW�9cV�9�W�9�X�9jW�9#V�9�W�9�V�9�U�9:X�9.Y�9�U�9�Y�9�[�9�V�9x   x   �T�9�S�9cW�9W�9T�98U�9�W�9�X�9Y�9�W�9W�9�X�9�Z�9eW�9�U�9�X�9�V�9�W�9�W�9�W�9�W�9hV�9�W�9�Y�91Y�9�V�9�V�9�Y�9>Z�9qX�9x   x   �V�9�V�9Z�9�V�9JV�9�W�92[�9�V�9�U�9bV�9V�9W�97X�9W�9�V�9�W�9�W�9�\�9�V�9�W�9W�9�V�9�X�9SW�9�U�9�V�9QV�9V�9_Y�9*X�9x   x   bW�9�X�9}Y�9�W�9�X�9�U�9�T�9�V�99Z�9�Y�9�X�9�U�9{V�9�X�9�W�9S�9EW�9RX�9PS�9�X�9�X�9�U�9�U�97X�9�Y�9�Y�9V�9�U�9�V�9KX�9x   x   �U�9YR�9�T�9�R�9W�9�W�9�Y�9wY�9�[�9�X�9�W�9CW�9U�9�W�9�Y�9�V�9GU�9�V�9FY�9�V�9cV�9JW�96X�9Y�9�[�9;Z�9\Y�9�V�9�V�9'S�9x   x   �V�9�V�9�V�9�R�9�W�9�W�9�X�9�V�9xT�9WS�9�W�9mX�9KW�9�W�9[�9Z�9]Y�9�[�9+Y�9W�9vW�9�W�9�R�9�T�9�V�9qX�9*X�9JX�9)S�9�U�9x   x   }x�9~��9���9��9܄�9M��9���9��9���9��9Y��9���9��9��9ρ�9H��9���9���9��9#��9Ä�9���9ց�9~��9u��9#��9���9�~�92��9�9x   x   |��9k��9t��9��9���9o�9���9��9`��9��9���9���9�}�9Ҁ�9��9���9���9~�9��9��9���9]��9��9��9��9���9|��9%�9z��9���9x   x   ���9t��9���9��9��9T��9v�9���9���9^~�9���9��9���9��9f~�9k��9E��9]��9��98�9i��9��9[�9ރ�9i��9*�9��9=��9]��9	��9x   x   ��9��9��9q}�9D��9���9X��9.��9��9Ԃ�9��9���9���9~��9���9���9X��9/��9Q��9`��9��9%��94��9���9b�9A�9��9��9>��9)��9x   x   ߄�9���9��9E��9���9e��9�9x��9��9A��9���9^��9���9���9��9��9R��9Ȃ�9���9���9=��9S��9���9Z��9���9E��96��9��9���9~�9x   x   J��9o�9U��9���9i��9��9"��9���9S��9���9X��9x��9ʂ�9���9:��9W��9���9k��9���9Ձ�9=��9r��9&��9��9��9ă�93��9v��9.��9ށ�9x   x   ���9���9y�9V��9���9'��9��9���94��9b��9���9^��9�9`��9���9���9��9ك�9 ��98��9��9��9��9k��9>��9���9���9	��9΂�9o��9x   x   ��9��9���9*��9s��9���9���9C��9���9̃�9���9��9;��9��9���9���9B��9���9��9��9���9���9�~�9Z��9	��92~�9���9��9�~�9g��9x   x   ���9c��9���9��9��9U��99��9��9΃�9���9��9̈́�9R��9���9*��9{��9��9���9���9���9��9���9��9���9=~�9�~�9��9m�9�~�9���9x   x   ��9��9^~�9ӂ�9=��9���9b��9˃�9���9���9[��9���9W��9���9��9)��9Y��9���9'��9�~�9��94��9���9Y��9W��9��9���9�~�9���95��9x   x   W��9���9���9��9��9S��9���9���9	��9^��9p��9Z��9���9��9Ȃ�9؆�9S��9P��9l��9���9��9��9_��9���9F��9���92��9"��9)��9L��9x   x   ���9��9��9���9^��9x��9_��9��9Ȅ�9���9Z��9���9#��9@��9��9���9���91��9��9ς�9/��9���9g��9���9��9��9S��9Q��9��9ƃ�9x   x   ��9�}�9���9���9���9Ȃ�9Ć�9?��9R��9Z��9���9&��9���9���9���9U��9��9�~�9���9{��9a��9���9��9��9ڄ�9S��9���9a��99��9Ղ�9x   x   ��9Ҁ�9��9|��9���9���9`��9��9���9���9��9A��9���9���9j��9\��90��9���9 ��9��9·�9��9Ä�9��9a��9���9ք�9=��9��9��9x   x   ΁�9��9e~�9���9��98��9���9~��9)��9��9Ƃ�9���9���9j��9�~�9���9��9̀�9��9m��9��9��9s��9���94��9.��9ԁ�9^��9ʀ�9��9x   x   E��9���9l��9���9��9V��9���9���9}��9,��9݆�9���9T��9Y��9���9%��9��9<��9^��9���9�9x��9��9@��97��9̃�9p��9 ��9C��9���9x   x   ���9���9D��9X��9S��9���9��9C��9��9V��9W��9���9��90��9��9��9A��9օ�9���9K��9���9���95��9���9���9t��9���9���9��9��9x   x   ���9
~�9^��9+��9�9h��9؃�9���9���9���9N��9.��9�~�9���9ʀ�9;��9ԅ�9�|�9ځ�9V��9ց�9���9Æ�9���9Ƀ�9(��9E~�9s��9���9ۀ�9x   x   ݅�9��9!��9R��9���9Ä�9��9��9���9)��9q��9���9���9���9��9_��9���9ځ�9e��9ԃ�9���9`��9���9$��9��9���9j��9���9��9��9x   x    ��9���9;�9_��9���9ׁ�9;��9	��9���9 �9���9Ђ�9{��9��9r��9���9M��9W��9҃�9���9F��9Ȃ�9���9���9��9���9��9Ё�9��9+��9x   x   �9���9j��9��9?��9;��9��9ƅ�9��9��9��92��9c��9ˇ�9��9Ä�9���9ԁ�9���9I��9���9C��9��9[��9��9^��9'��9��9���9ς�9x   x   ���9Y��9
��9"��9X��9t��9��9���9���94��9��9���9���9��9��9x��9���9���9`��9Ȃ�9>��94��9'��9j��9��9׃�9��9!��9k��9c��9x   x   ҁ�9��9]�9/��9���9"��9��9�~�9��9���9d��9g��9
��9���9m��9��9;��9Æ�9���9���9��9)��9N��9���9T��9W��9��9���9j��9E��9x   x   |��9��9��9���9U��9��9g��9]��9���9X��9���9��9��9��9���9<��9���9���9"��9���9]��9l��9���9+��9$��9���9��9Ԅ�9w��9Æ�9x   x   v��9��9k��9^�9�9��9?��9��9=~�9]��9G��9 ��9݄�9a��94��97��9���9Ƀ�9���9���9��9��9U��9&��9<��9ʂ�9��9��9�|�95��9x   x   !��9���9)�9C�9B��9Ã�9���9/~�9�~�9���9���9��9V��9���9+��9̓�9w��9)��9���9���9^��9؃�9U��9���9ɂ�9���9*��9}��9!~�9���9x   x   ���9z��9��9��98��96��9���9���9��9���92��9P��9���9ׄ�9ҁ�9s��9���9B~�9k��9��9%��9��9��9��9��9+��9��9���9q��9���9x   x   �~�9&�9?��9��9��9{��9	��9��9l�9�~�9%��9M��9^��98��9c��9��9���9w��9���9Ӂ�9��9 ��9���9҄�9��9}��9���9���9'��9��9x   x   /��9t��9X��9:��9���9.��9΂�9�~�9�~�9���9'��9��9=��9��9π�9C��9��9���9��9��9���9k��9g��9u��9�|�9!~�9r��9$��9��9��9x   x   ˂�9���9��9-��9~�9��9m��9d��9���97��9N��9ȃ�9Ղ�9���9~��9���9���9ڀ�9��9+��9ς�9a��9E��9�92��9���9���9��9��9΅�9x   x   ���9���9���9M��9x��9\��96��9)��9°�9��9���9���9���9��9���90��9J��94��9.��9W��9���9s��9I��9��9���9o��9;��9а�9|��9���9x   x   ���9X��9���9@��9M��9p��9���9���9���9���9���9)��9��9^��9|��9ϰ�9���9n��9ݮ�9-��9���9���9��9E��9<��9���9��9��9E��9���9x   x   ���9���9��9���9s��9j��9���9��9���9���9گ�9���9��90��9���9X��9&��9w��9���9��9խ�9���9z��9���9���9Y��9���9Į�9g��9]��9x   x   M��9?��9���9��9*��9 ��9	��9G��9ڮ�9���9���9���9���97��9y��9]��9j��9D��9t��9��9���9���9��9���9_��9{��9׭�9T��9	��9��9x   x   x��9M��9p��9.��9M��9G��9���9w��9���9���9���9p��9ܬ�9���9D��9V��9���9���9���9Q��9���9®�97��9��9-��9L��9]��9z��9u��9\��9x   x   _��9p��9h��9���9F��9���9ư�9���9��9.��9���9���9���9��90��9̰�9R��9��9��9���9���9"��9Ʈ�9#��9r��9��9��9]��9O��9$��9x   x   5��9���9���9��9���9ʰ�9���9o��9ݯ�9c��9W��9F��9���9��9~��9��9F��9{��9ٯ�9��9���9���9���9t��9v��9/��9���9���9N��9��9x   x   -��9���9��9L��9w��9���9k��9���9֮�9A��9��9��9:��9���9!��9ڮ�9֯�9ׯ�9���9���9���9��9��9���9Q��9ݳ�9���9��9���9c��9x   x   ɰ�9���9��9׮�9���9��9گ�9׮�9r��9���9��9 ��9���9��9ܫ�9E��9 ��9��9��9ծ�9���9��9��9��9���9���9���9I��9��9��9x   x   ��9���9���9���9���9,��9e��9>��9���9���9f��9���9���9-��9��9r��9���9-��9P��9;��9o��9
��9��9��9A��9H��9p��9i��9��9��9x   x   ���9���9ׯ�9���9���9���9U��9
��9��9h��9��9U��9��9���9���9��9ʬ�96��9>��9��9��9���9���9q��9��9��9��9M��9@��9M��9x   x   ���9)��9���9���9u��9���9D��9��9 ��9���9Y��9���9O��9��9B��9	��9���9���9B��9ڮ�9C��9?��9���9���9<��93��9��9~��9=��9��9x   x   ���9��9��9���9ܬ�9���9���98��9���9���9 ��9L��9I��9��9ū�9 ��9ɰ�9M��9U��9���9���9>��9��9���9���9���9��9��9��9���9x   x   ��9]��92��97��9���9��9��9���9��9+��9���9��9��9\��9���9��9H��9���9ɯ�9���9���9���9��9���9ݰ�9���9��9 ��9��9���9x   x   ���9}��9���9z��9B��90��9}��9#��9��9��9���9B��9ƫ�9���9z��9��9��9c��91��9˱�9���9��9ˮ�9p��9��9���9��9P��9F��9$��9x   x   4��9Ͱ�9X��9^��9X��9Ͱ�9��9ٮ�9D��9s��9��9��9��9޳�9��9j��9���9ͱ�9L��9���9��9���9y��9s��9��9���9��9��9���9���9x   x   Q��9���9&��9j��9���9S��9E��9ׯ�9 ��9 ��9Ǭ�9���9̰�9E��9��9���9l��9K��9���9ܭ�9���9���9ΰ�9,��9j��9��9��9���9��9ί�9x   x   4��9m��9z��9@��9���9��9y��9گ�9��9+��92��9���9O��9���9d��9ͱ�9R��9S��9J��9��9D��9��9���9���92��9���9��9I��9:��9Į�9x   x   -��9ޮ�9���9v��9î�9���9ԯ�9���9��9S��9>��9E��9T��9˯�90��9E��9���9F��9q��99��9*��9���9��9���9���9���9��9L��9F��9���9x   x   Y��9*��9��9��9M��9���9��9���9ծ�9=��9	��9ޮ�9���9���9̱�9���9߭�9��99��9��9���9���9���9���9��9O��9���9��9i��9S��9x   x   ���9���9֭�9���9���9���9���9{��9���9w��9��9B��9���9���9���9��9���9F��9-��9���9-��9���9\��9ұ�9^��9���9U��9���9��9���9x   x   s��9���9���9���9���9#��9���9��9��9��9���9;��9<��9���9��9���9���9��9���9���9���9Ү�9N��9���9��97��9���94��9���9:��9x   x   L��9
��9z��9��96��9Ʈ�9���9��9	��9��9���9���9 ��9��9ή�9{��9ΰ�9���9��9���9\��9L��9��9��9���9h��9B��9>��9���9���9x   x   	��9G��9���9���9��9&��9s��9���9��9��9m��9 ��9���9���9p��9n��9+��9���9���9���9ұ�9���9��9���9e��9@��9���9;��9���9���9x   x   ��99��9���9c��9/��9s��9t��9O��9��9A��9���9C��9��9װ�9��9��9j��94��9���9 ��9^��9 ��9���9e��9���9ŭ�9b��9?��9��9���9x   x   u��9���9W��9{��9I��9��91��9��9���9I��9��94��9���9���9���9���9��9���9���9N��9���9;��9i��9=��9���9���9���9��9���9���9x   x   9��9��9���9֭�9^��9��9���9���9���9r��9{��9��9��9��9���9��9��9��9���9���9X��9���9A��9���9a��9���9 ��9߯�9	��9���9x   x   Ұ�9���9Ʈ�9S��9x��9\��9���9��9F��9j��9R��9���9ۭ�9��9O��9��9���9B��9K��9��9���95��9B��9>��9E��9��9ܯ�9\��93��9���9x   x   ��9B��9l��9��9t��9O��9M��9���9��9��9=��9?��9��9��9F��9��9��9:��9G��9e��9��9���9���9���9��9���9��94��9��9��9x   x   ���9���9]��9��9\��9%��9��9f��9	��9��9J��9	��9���9���9*��9��9ү�9Ȯ�9���9O��9���9:��9���9���9���9���9���9���9��9y��9x   x   ���93��9���9U��9���9r��9u��9b��9)��9���9}��9��9���9l��9���9>��9m��9���9���94��9��9���9
��9���9d��9���9���9$��9���9|��9x   x   .��9e��9���9)��9���9���9<��9x��9���9o��9l��9���9��9��9���9���9���9���9F��9���9E��9���9��9���9L��9 ��9I��9���9��9���9x   x   ���9���9*��9���9I��9o��9��9���9���9"��9���90��9���9���9Y��9
��9���9���96��9m��9t��9��9���9���9���9w��9���9���9��9��9x   x   U��9,��9���9��9e��9���9���99��9*��9T��9��9'��9���9\��9?��9���9���9���9���9���9A��9���9���9���9���9��9b��9���9Z��9h��9x   x   ���9���9I��9g��9x��9���9���9���9���9���9M��9���9"��9x��99��98��9���9���9���9���9���9O��9g��9���9Y��9���9���9,��9m��9���9x   x   q��9���9l��9���9���9b��9y��9���9���9��96��9���9s��9M��9���9@��9)��9r��9x��9}��9D��9y��9��9���9���9O��9��9G��9V��9 ��9x   x   s��9=��9��9���9���9u��9b��9��9��9l��9?��9���9��9���9���9���98��9���9��9���9���9��9d��9��9���9^��9���9���9��9c��9x   x   a��9u��9���9>��9���9���9��9��94��9���93��95��9$��9N��9���9��9 ��9	��9���9���9n��9)��9��9���9���9���9(��9���9���9v��9x   x   *��9���9���9)��9���9���9 ��98��9���9p��9���9���9��9���9h��9���96��9���9���9z��9{��9��9J��9D��9C��9u��9*��9��9?��9��9x   x   ���9s��9*��9W��9���9��9m��9���9r��9���9���9���9���9���9���9���9C��9���9���9V��9���9���9���9���9r��9E��9%��9���9%��9���9x   x   {��9j��9���9��9I��93��9B��91��9���9���9���9d��9��9���9���9��9|��9���95��9/��9R��9���9��9���9���9��9E��9@��9o��9���9x   x   ��9���9.��9&��9���9���9���98��9���9���9f��9=��9O��9	��9���9��9���9���9��9��9���9���95��9���9n��9���9k��9���90��9q��9x   x   ���9!��9���9���9!��9q��9��9&��9
��9���9��9O��9D��9��9���9���9���9���9P��9"��9��9���9x��9v��9?��9*��9���9���9��90��9x   x   m��9��9���9Z��9w��9L��9���9O��9���9���9���9	��9��9/��9��9���9F��9��9D��9'��9]��9���9���9��9���9L��9���9b��9���9M��9x   x   ���9���9Y��9>��94��9���9���9���9d��9���9���9���9���9��9;��9���9k��9 ��9o��9F��9���9v��9���9���9{��9A��9���9|��9���9Q��9x   x   <��9���9��9���98��9=��9���9��9}��9���9��9��9��9���9���9���9���9V��9z��9I��9��9���90��9��9���9?��9���9��9���9w��9x   x   m��9���9���9���9���9(��98��9���95��9G��9���9���9���9F��9i��9���9���9Y��9���9.��9���9@��9���9<��9���9q��9���9%��95��9S��9x   x   ���9���9���9���9���9s��9���9
��9���9���9���9���9���9��9��9T��9]��9���9���9��9���9���9���9���9R��9���9M��9���9���99��9x   x   ���9E��94��9���9���9v��9��9���9���9���94��9��9M��9H��9p��9z��9���9���9���9���9��9w��9W��9A��9���9���9S��9��91��9���9x   x   7��9���9l��9���9���9���9���9���9}��9O��9.��9��9 ��9#��9D��9J��9/��9��9���9���9u��9���9?��9���9[��9u��9���9���9���97��9x   x   ��9G��9s��9H��9���9E��9���9q��9{��9���9O��9���9	��9\��9���9��9���9���9��9n��9���9���9��9���9���9��9Y��9���9i��9%��9x   x   ���9���9��9���9N��9x��9
��9!��9���9���9���9���9���9���9v��9���9;��9���9|��9���9���9���9j��9���9��9���9��9���9���9
��9x   x   
��9��9���9���9g��9��9a��9��9K��9���9��98��9u��9���9���90��9���9���9U��9=��9��9h��9t��9���9���9~��9���9���9��9���9x   x   ���9���9���9���9���9���9��9���9G��9���9���9���9t��9
��9���9���9=��9���9A��9���9���9���9���9E��9���9_��9;��9���9���9���9x   x   d��9M��9���9���9S��9���9���9���9C��9t��9���9i��9<��9���9|��9���9���9P��9���9Z��9���9��9���9���9���9}��9���9���9���9���9x   x   ���9��9z��9��9���9O��9_��9���9u��9H��9��9���9.��9J��9:��9A��9o��9���9���9r��9��9���9~��9c��9���9K��9���98��9���9��9x   x   ���9M��9���9b��9���9��9���9(��9+��9&��9F��9i��9|��9���9���9���9���9L��9R��9���9V��9��9���9=��9���9���9���9K��9��9��9x   x   ��9���9���9���9,��9K��9���9���9��9���9?��9���9���9f��9~��9��9(��9���9��9���9���9���9���9���9���97��9I��9��9���9���9x   x   ���9��9��9[��9m��9Z��9��9���9B��9$��9l��94��9��9���9���9���92��9���9.��9���9i��9���9��9���9���9���9��9���9���9��9x   x   y��9���9��9e��9���9 ��9a��9r��9��9���9���9q��96��9Q��9M��9w��9V��97��9���9>��9'��9��9���9���9���9��9��9���9��9��9x   x   ��9��9	�9	�9��9��9f
�90�9�9	�9��9:�9��9��9��9��9:�9��9��9��9��9L�9<�9��9��9W�9��9��9w	�9�9x   x   ��9��91�9��9	�97�9�
�9��9�9B
�9��9��9w�9��94�9��9��9�98�9-�9d�9��9�
�9�9�	�9�9��9+�9V�9.�9x   x   	�91�9�	�9�
�9Q
�9��9V�9��9��9�
�9��9��9~�9t�9��9��9�9��9<�9�
�9��9%�9��9��9A�9�
�9�	�9��9�9h�9x   x   	�9��9�
�9>�9r�9��9��9�9.�9��9x�9�92�9��9��9��9 
�9*�9��9�	�9�9��9v�9��9��9��9c�9�	�9��9��9x   x   ��9�9O
�9t�9"�9t�9!�98�9��9��9;
�9��9I�9+�9��9t�9H�94�9o�9��9�
�9��9��9u�9
�9��9g�9��9��9��9x   x   ��9:�9��9��9~�91�9��9��90�9�99�9��9{�9��9,�9�9�9[�9�9��9f�9��9��9��9�	�9�9��9O�9��9��9x   x   b
�9�
�9Y�9��9!�9��9k
�9Z�93
�9p�9��9Q�9��9��9~�9T�9��9�9`	�9E�9��9��9�
�9��9�
�9�
�9M�9#�9��9�
�9x   x   .�9��9��9�9<�9��9Z�9l�9u
�9��9.�9��9a�9��9)�9
�9�
�9u�9:�9f�9��9q�9|	�9��9��9>�9Y�9��9o�9�9x   x   �9�9��9/�9��93�93
�9r
�9z�96�9}�9s�9��9u
�9	�9�
�9C
�96�9��9��9	�9U�9��92�9��9�9��9J�9!�9��9x   x   �9C
�9�
�9��9��9	�9m�9��98�9x�9|�9i�9��9�
�98�9��9�9��9{�9[�9�9��9�
�9��9��9��9F�9+�9��9�	�9x   x   ��9��9��9y�9>
�9=�9��9)�9}�9��9F�9f�9��9��9X�9��9�	�9��9;�9Q�98�9(�9�9��94�9�
�9C�9�9H�9��9x   x   ?�9��9��9�9��9��9R�9��9t�9h�9c�9S�9}�9�9��9��9-	�9,�9��9��9��9�9��9o�9��9��9��9��9v�9#�9x   x   ��9s�9~�93�9N�9{�9��9\�9��9��9��9~�9��9
�9��9��9��9m�9u�9p�9)�9��9n�9w�9��9��9��9�9U�9@�9x   x   ��9��9v�9��9.�9��9��9��9x
�9�
�9��9�9�99�9��9�9��96�9��9��94�9��9%�9f�9.�9^�9�9��9j�9�9x   x   ��99�9��9��9��9*�9{�9'�9�99�9T�9��9��9��9��9��9F�9��9�9��9�	�9!�9T�9-�9��9��9�	�9T�9A�9��9x   x   ��9��9��9��9{�9�9T�9
�9�
�9��9��9��9��9�9��9��96�9��9�9��9v�9�9�92�9|�9��9�9<�9��9�9x   x   6�9��9�9
�9I�9�9��9�
�9B
�9�9�	�9+	�9��9��9E�9:�9P�9��9��9��9��9��9\�9��9_�9�9��9��9�9��9x   x   ��9�9��9)�9.�9`�9�9u�94�9��9��9+�9q�96�9��9��9��9��9��9��9��9 �95�9��9��9�9��9�96�9}�9x   x   ��90�9?�9��9m�9�9]	�9>�9��9}�9@�9��9s�9��9�9�9��9��9��9��9�9�9t�9��9"�9��9��9d�9��9��9x   x   ��91�9�
�9�	�9��9��9A�9c�9��9]�9U�9��9q�9��9��9��9��9��9��9.�9Q�9��9��9E�9G�9w�9#�9+�95�9��9x   x   ��9a�9��9�9�
�9f�9��9��9	�9�98�9��9*�93�9�	�9x�9��9��9�9T�9��9t�9�9��9I�9��9�
�9m�9
�9��9x   x   K�9��9*�9��9��9��9��9u�9U�9��9/�9�9��9��9"�9�9��9�9�9��9n�9p
�9��9��9Y�9��9��9��9��9��9x   x   :�9�
�9��9w�9��9��9�
�9�	�9��9�
�9�9��9m�9$�9P�9	�9`�92�9r�9��9�9��9?�9%�9��9��9	�9��9D�9_�9x   x   ��9	�9��9��9u�9��9��9��92�9��9��9r�9w�9j�9,�92�9��9��9��9F�9��9��9%�9��9W�9t�9�9��9��9��9x   x   ��9�	�9D�9��9
�9�	�9�
�9��9��9��97�9��9��9,�9��9|�9[�9��9�9B�9D�9T�9��9Q�9�9��9��9��9��9u�9x   x   P�9��9}
�9��9��9��9�
�9;�9�9��9�
�9��9��9_�9��9��9!�9!�9��9{�9��9��9��9r�9��9��9�9[�9��9
�9x   x   ��9��9�	�9j�9g�9��9M�9X�9��9D�9F�9��9��9�9�	�9�9��9��9��9!�9�
�9��9
�9�9��9�9/�9>�9d�9��9x   x   ��9-�9��9�	�9��9O�9$�9��9M�9+�9�9��9�9��9W�9>�9��9�9d�9*�9m�9��9��9��9��9^�9?�93
�9��9<�9x   x   u	�9W�9�9��9��9��9��9o�9#�9��9I�9u�9R�9e�9E�9��9�97�9��92�9�9��9I�9��9��9��9f�9��9p�9��9x   x   �90�9c�9��9��9��9�
�9�9��9�	�9��9#�9@�9�9��9�9��9~�9��9��9��9��9]�9��9q�9
�9��9<�9��9$�9x   x   �B�9^?�9J>�9�@�9~9�9�?�9�=�9�<�9�>�9�?�9�@�9s<�9K@�9jA�9�=�9I>�9�=�9�B�9@�9�=�9@�9�>�9{>�9)<�9P>�9�?�9:�9�@�9�=�9V?�9x   x   \?�9�>�9�?�9�=�9�;�9�>�9�A�9�=�9�;�9F=�9)B�9b:�9?�9�>�9_;�9�<�9�=�9�=�9�:�9�A�9z>�9�;�9�>�9�A�9d>�9e;�9=�9�?�9c?�9�@�9x   x   N>�9�?�9@>�9�@�9�<�9�@�9P?�9�>�9g?�9~>�9a@�9�;�9�>�9U=�9b>�9 =�9@�9S<�9�?�9�>�9�>�9>�9#?�9�@�9n=�9�@�9�>�9(@�98<�9 7�9x   x   �@�9�=�9�@�9u>�9�=�9�<�9P<�9$>�9d>�9�=�9�<�9�?�9�=�9^?�9�>�9�=�9�>�9a<�9�>�9�=�9�?�9�<�9v<�9W=�9>�9�@�9q<�9�A�9/>�9�<�9x   x   �9�9�;�9�<�9�=�9�;�9�<�9�?�9�<�90A�9�?�9�>�9�A�9.>�91B�9�>�9�@�9�?�9�?�9!A�9�<�9T>�9�<�9<�99>�9�<�9U<�9)9�9<�9�<�9^=�9x   x   �?�9�>�9�@�9�<�9�<�9�@�9�?�9�<�9=A�9�?�9�?�9�:�9�>�9i>�9�:�9@@�9
?�9�@�9�=�9@�9;B�9U<�9�;�9%A�9>�9@�9M>�9F;�9;�9�=�9x   x   �=�9�A�9Q?�9N<�9�?�9�?�9n=�9�?�9�<�9�;�9�<�9&=�9�A�9�<�9�<�9�:�9q>�9s?�9�<�9P?�9�>�9�=�9�>�9jB�9�=�9c@�9?�9�<�9�>�99A�9x   x   �<�9�=�9 ?�9%>�9�<�9�<�9�?�9NE�9�A�9�>�9�A�9�<�9�=�9�A�9?�9vA�9D�9U@�9�=�9_=�9>�9�>�9�=�9�<�9t:�9A�9:�9�:�9	A�9�9�9x   x   �>�9�;�9h?�9f>�93A�98A�9�<�9�A�9jA�9^?�9C�9�>�9EB�9?�9tA�9hA�9�=�9o@�9�@�9�>�9b>�9%<�9v>�9�<�9Z@�9qA�97�9�@�9Z@�9�<�9x   x   �?�9E=�9|>�9�=�9�?�9�?�9�;�9�>�9_?�9=�9�>�9�>�9E>�9&?�9�>�9�;�9?�9�@�9�<�9A?�9>�9�>�9�>�9!=�9�>�9=<�9D<�9p?�9Q=�9�=�9x   x   �@�9,B�9b@�9�<�9�>�9�?�9�<�9�A�9C�9�>�9=�9�>�9@B�9�A�9
<�9�?�9�>�9f=�9z@�9�@�9�@�9p?�9
<�9�>�9�>�9RA�9N>�9�=�9�<�9n?�9x   x   t<�9c:�9�;�9�?�9�A�9�:�9%=�9�<�9�>�9�>�9�>�9�>�9�=�9A=�99;�9FB�9 >�9�;�9 ;�9n=�9x>�9d?�9T@�9�?�9�>�9?�9A�9]@�9C?�9>�9x   x   G@�9?�9�>�9�=�9,>�9�>�9�A�9�=�9DB�9A>�9=B�9�=�9{@�9&?�9�<�9?�9q@�9>�9�?�9�=�9�=�9:>�9�>�9�A�9�?�9t@�9�>�9�=�96>�9I?�9x   x   kA�9�>�9U=�9]?�90B�9j>�9�<�9�A�9?�9'?�9�A�9E=�9(?�9MC�9
?�9D;�9�>�9B�9�>�9?�9�?�9�<�9�?�9�>�9@�9H@�9�<�9c@�9^=�9�=�9x   x   �=�9^;�9d>�9�>�9�>�9�:�9�<�9!?�9nA�9�>�9<�98;�9�<�9?�9�?�9;<�9�=�9�=�97=�9BB�9�A�9�B�9U?�9�<�9e>�9PB�9YA�9?C�9Y>�9e>�9x   x   K>�9~<�9�<�9�=�9�@�9?@�9�:�9uA�9aA�9�;�9�?�9CB�9?�9B;�9;<�9y=�9�?�9{?�9?�9H>�9]A�9 >�96A�9�@�9�>�9XB�9W=�9o>�9^>�9f?�9x   x   �=�9�=�9@�9�>�9�?�9
?�9j>�9D�9�=�9?�9�>�9>�9r@�9�>�9�=�9�?�9�?�9?�9�=�9�>�9�>�91=�9�>�9>�9"=�9)?�9�>�9�?�9�@�9�>�9x   x   �B�9�=�9Y<�9a<�9�?�9�@�9s?�9X@�9r@�9�@�9d=�9�;�9>�9B�9�=�9|?�9?�9�A�9D�9y=�9B�9�@�9v?�9ZB�9
>�9]C�9aA�9{>�9�?�9�=�9x   x   @�9�:�9�?�9�>�9"A�9�=�9�<�9�=�9�@�9�<�9w@�9;�9�?�9�>�93=�9?�9�=�9 D�9�?�9�=�9C�9�>�9OC�9g>�9�?�9�D�9�>�9�>�9�=�9�=�9x   x   �=�9�A�9�>�9�=�9�<�9@�9P?�9^=�9�>�9A?�9�@�9p=�9�=�9?�9?B�9H>�9�>�9v=�9�=�9�D�9�A�9�B�9[C�9=�9]>�9�=�9�>�9=B�9 ?�9�=�9x   x   @�9|>�9�>�9�?�9X>�9@B�9�>�9>�9c>�9>�9�@�9t>�9�=�9�?�9�A�9\A�9�>�9B�9C�9�A�9�@�9�A�9E�9�A�9�>�9aA�9�A�9v?�9q>�9>�9x   x   �>�9�;�9>�9�<�9�<�9X<�9�=�9�>�9&<�9�>�9o?�9_?�9:>�9�<�9�B�9>�90=�9�@�9�>�9�B�9�A�9�=�9�?�9�<�9?�9:B�9%=�9>�9�>�9�@�9x   x   z>�9�>�9"?�9s<�9 <�9�;�9�>�9�=�9v>�9�>�9<�9U@�9�>�9�?�9W?�93A�9�>�9w?�9NC�9_C�9E�9�?�97@�93@�9�>�9�?�9�>�9�@�9�;�9�>�9x   x   ,<�9�A�9�@�9W=�97>�9#A�9eB�9�<�9�<�9!=�9�>�9�?�9�A�9�>�9�<�9�@�9>�9`B�9h>�9=�9�A�9=�95@�9�=�9	?�9�A�9/@�9W?�9g<�97=�9x   x   R>�9c>�9p=�9>�9�<�9>�9�=�9v:�9[@�9�>�9�>�9�>�9�?�9@�9h>�9�>�9=�9
>�9~?�9^>�9�>�9?�9�>�9?�9�?�9?�9q=�9p?�9�@�9�9�9x   x   �?�9e;�9�@�9�@�9S<�9@�9d@�9A�9rA�9=<�9TA�9?�9v@�9F@�9PB�9WB�9)?�9]C�9�D�9�=�9aA�9;B�9�?�9�A�9?�9(B�9E<�9�@�9�@�9�@�9x   x    :�9=�9�>�9o<�9)9�9R>�9?�9:�97�9G<�9N>�9A�9�>�9�<�9VA�9W=�9�>�9`A�9�>�9�>�9�A�9!=�9�>�94@�9q=�9G<�977�9�:�9`?�94=�9x   x   �@�9�?�9'@�9�A�9<�9D;�9�<�9�:�9�@�9n?�9�=�9]@�9�=�9e@�9?C�9l>�9�?�9z>�9�>�9@B�9x?�9>�9�@�9W?�9o?�9�@�9�:�9�;�9�;�9�<�9x   x   �=�9^?�9:<�94>�9�<�9;�9�>�9
A�9^@�9O=�9�<�9A?�9:>�9`=�9X>�9[>�9�@�9�?�9�=�9!?�9r>�9�>�9�;�9h<�9�@�9�@�9\?�9�;�9x<�9�=�9x   x   V?�9�@�97�9�<�9c=�9�=�98A�9�9�9�<�9�=�9l?�9>�9K?�9�=�9i>�9h?�9�>�9�=�9�=�9�=�9	>�9�@�9�>�98=�9�9�9�@�91=�9�<�9�=�9S7�9x   x   i�9�l�9jr�9�p�9p�9�q�9*q�9�n�9kq�9[q�9�o�9�q�9�q�9�o�9ms�9hq�9�r�9p�9zr�9%r�9�o�9rp�9�q�9^o�9q�9�p�9�p�9~q�9�q�9�l�9x   x   �l�9}j�9Km�9]l�9]o�9�n�9�m�9�s�9\q�9r�9�p�9�t�95t�9�o�9t�9u�9�o�9ts�9�t�9�o�9�r�9�r�9�r�9�m�9ro�9*o�9�k�91m�9:k�9�l�9x   x   er�9Gm�9�m�9*o�9�q�9�k�9�m�9fm�9p�9np�9�l�9xs�9�o�9�p�9v�9p�9Vp�9�s�9+m�9�p�9�n�9;m�9�n�9�k�9�q�9vo�9�m�9Sm�91q�9t�9x   x   �p�9^l�9,o�9;n�9�n�95r�9�r�9�o�9Ot�9�p�9�r�9dt�9an�9�p�9rp�9�n�9Lt�9�q�9=p�9�t�9�p�9�r�9�q�9�n�9>n�9!o�9�k�9�q�9�q�95p�9x   x   p�9[o�9�q�9�n�9�s�9#s�9eq�98q�9
o�9�o�9�p�9�r�9�r�9p�9�r�9�q�9bq�9mp�9bn�94q�9%q�9�r�9�t�9io�9Nq�9�o�9<p�9�o�9?j�9�q�9x   x   �q�9�n�9�k�97r�9s�9Vg�9.p�9�o�9�n�9�q�9an�9�r�9�o�9go�9os�9�n�9�p�90o�9�o�9�o�9Gh�9s�9�p�9l�9�n�9q�9q�9�r�9<r�9p�9x   x   *q�9�m�9�m�9�r�9dq�9.p�9�u�9�l�9pq�9�r�9�r�9}r�94q�9\r�9�r�9�r�9�q�9il�9~v�9p�9xp�9}s�9�n�9�m�9Oq�9Dn�9`l�9qx�9�l�9�n�9x   x   �n�9�s�9bm�9�o�93q�9�o�9�l�9hm�9wo�9�n�9�o�9tp�9$q�9�o�9�n�9p�9�l�9�l�9^o�9�q�93p�9�l�9�r�9�n�9�q�9m�9Rq�9�q�9�l�9sp�9x   x   mq�9Zq�9p�9Lt�9o�9�n�9sq�9vo�9Do�9�p�9o�9+r�9bn�9*q�9�n�9o�9�r�9�n�9�n�9�t�9�o�9�q�9�r�9�o�9�n�94r�9^t�9/q�9@o�9	q�9x   x   Yq�9 r�9qp�9�p�9�o�9�q�9�r�9�n�9�p�9Gm�9�q�9�q�9�m�9�p�9�o�9cr�9�p�9�p�9�o�9np�9�r�9p�9vt�9's�9�n�9�o�9�p�9ao�96r�9/t�9x   x   �o�9�p�9�l�9�r�9�p�9`n�9�r�9�o�9o�9q�9u�9�q�9�n�9o�9dr�9!o�9�p�9~r�9@m�9p�9-p�9�n�9q�9/q�9�q�9�t�9q�9�p�9�q�9�n�9x   x   �q�9�t�9ws�9et�9�r�9�r�9|r�9tp�9(r�9�q�9�q�9=r�9	q�9�r�9s�9r�9�s�9�s�9�t�9hq�9jq�9�r�9�p�9�l�9�o�9p�9�m�9sq�9r�9�p�9x   x   �q�96t�9�o�9fn�9�r�9�o�9/q�9#q�9en�9�m�9�n�9	q�9mp�9�o�9Xr�9Ko�9�p�9�s�9�r�9(q�9r�9�q�9�r�9p�9q�9o�9�q�9Tq�9Ns�9
r�9x   x   �o�9�o�9�p�9�p�9p�9jo�9Vr�9�o�9*q�9�p�9}o�9�r�9�o�9_p�9[p�9to�9p�9!o�9�n�9�s�9�o�9�q�9�q�9jp�9\q�9�r�9�r�9�o�9�q�93o�9x   x   qs�9
t�9v�9tp�9�r�9qs�9�r�9�n�9�n�9�o�9er�9s�9Xr�9Zp�9�v�9�t�9�s�9ns�9Aq�9�q�9tq�9�q�9o�9u�9n�9�p�9�p�9er�9�q�9�s�9x   x   hq�9u�9p�9�n�9�q�9�n�9�r�9p�9o�9ar�9!o�9r�9Ko�9xo�9�t�9Ip�9�r�9tr�9�p�9.q�9�q�9Hn�9�v�9�v�9]o�9�r�9�p�9�p�9uq�9kr�9x   x   �r�9�o�9Wp�9Nt�9aq�9�p�9�q�9�l�9�r�9�p�9�p�9�s�9}p�9p�9�s�9�r�9�o�9r�9�r�9s�9Nt�9�r�9yo�99s�9�r�9qs�9�r�9�q�9q�9�r�9x   x   p�9ps�9�s�9�q�9lp�90o�9kl�9�l�9�n�9�p�9~r�9�s�9�s�9 o�9ps�9sr�9!r�9?s�9o�9�o�9u�9q�9Pp�9Lu�9rp�9,o�9�s�9�q�9�q�9�s�9x   x   zr�9�t�9*m�9@p�9]n�9�o�9�v�9Xo�9�n�9�o�9Bm�9�t�9�r�9�n�9Cq�9�p�9�r�9o�9�p�9�s�9�o�9�t�98p�9~t�9�o�9�n�9s�9�p�9r�9}n�9x   x   #r�9�o�9�p�9�t�92q�9�o�9p�9�q�9�t�9mp�9p�9jq�9"q�9�s�9�q�90q�9s�9�o�9�s�9_m�9�o�9Fp�9.l�9�s�9[q�9�r�9Bq�9�q�9�r�99q�9x   x   �o�9�r�9�n�9�p�9&q�9>h�9yp�97p�9�o�9�r�9.p�9mq�9r�9�o�9yq�9�q�9Qt�9u�9�o�9�o�9�n�9�o�9Kq�9�t�9Js�9or�9	q�9�o�9Ts�9�p�9x   x   qp�9�r�96m�9�r�9�r�9s�9{s�9�l�9�q�9p�9�n�9�r�9�q�9�q�9�q�9En�9�r�9q�9�t�9Gp�9�o�9)t�9Lp�9ls�9o�9�p�9�r�9�q�9�q�9*o�9x   x   �q�9�r�9�n�9�q�9�t�9�p�9�n�9�r�9�r�9tt�9q�9�p�9�r�9�q�9o�9�v�9zo�9Pp�96p�9,l�9Kq�9Jp�9p�9>v�9�n�9r�9#r�9q�9r�9t�9x   x   co�9�m�9�k�9�n�9go�9l�9�m�9�n�9�o�9)s�9.q�9�l�9p�9hp�9	u�9�v�9:s�9Gu�9{t�9�s�9�t�9ks�9>v�9�u�9�p�9�o�9[m�9�p�9�q�9Aq�9x   x   
q�9oo�9�q�9;n�9Mq�9�n�9Oq�9�q�9�n�9�n�9�q�9�o�9q�9_q�9n�9_o�9�r�9wp�9�o�9^q�9Ls�9o�9�n�9�p�9�p�9p�9�p�9�o�9o�94p�9x   x   �p�9.o�9|o�9$o�9�o�9q�9An�9m�90r�9�o�9�t�9p�9#o�9�r�9�p�9�r�9ns�9&o�9�n�9�r�9kr�9�p�9�q�9�o�9p�9�t�9�p�9tq�9�l�9`o�9x   x   �p�9�k�9�m�9�k�9?p�9q�9[l�9Rq�9\t�9�p�9q�9�m�9�q�9�r�9�p�9�p�9�r�9�s�9!s�9Bq�9q�9�r�9r�9am�9�p�9�p�9�s�9-r�9hl�9:p�9x   x   |q�9.m�9Um�9�q�9�o�9s�9rx�9�q�9/q�9ao�9�p�9uq�9Rq�9�o�9dr�9�p�9�q�9�q�9�p�9�q�9�o�9�q�9q�9�p�9�o�9wq�92r�9�w�9s�9Gp�9x   x   �q�9=k�94q�9�q�9Aj�9>r�9�l�9�l�9=o�94r�9�q�9!r�9Ms�9�q�9�q�9sq�9q�9�q�9 r�9�r�9Qs�9�q�9r�9�q�9o�9�l�9jl�9s�9qj�9�p�9x   x   �l�9�l�9 t�90p�9�q�9p�9�n�9qp�9q�90t�9�n�9�p�9r�93o�9�s�9ir�9�r�9�s�9{n�9>q�9�p�9+o�9t�9Cq�96p�9bo�9?p�9Bp�9�p�9�t�9x   x   ��9���9L��9 ��9̥�9���9��9���9r��9ۡ�9q��9s��9���9��9���9��9p��9���9���9���9[��9v��9h��9_��9���9a��9i��9���9I��9v��9x   x   ���9���9��9��9;��9��9G��9��9��9���9���9��9#��9��9���9���9C��9M��9��9���9a��9��9I��9���9��9;��9y��9��9r��9��9x   x   M��9��9٧�9e��9��9���9���9ƥ�9ģ�9���9k��91��9"��9ب�9;��9/��9"��9:��9��9#��9'��9���9#��9��9���9���9��9���91��9L��9x   x    ��9��9b��9w��9��9���9��9���9��9���9p��9R��9��9Ӥ�9Q��9���9-��9k��9���9���9h��9Z��9¢�9"��9���9)��9)��9Ɯ�9���9���9x   x   ̥�9>��9��9��9ʞ�9���9ʤ�9���9<��9��9W��9n��9���98��9��9���9s��9��9a��9���9c��9@��98��9��9ե�95��9w��9#��9#��9
��9x   x   ���9���9���9���9���95��9��9u��9զ�9=��9M��9��9���9��9ƥ�9r��9���9���9d��9 ��9���9��9G��9s��9���9���9���9n��9���9���9x   x   ��9H��9���9��9ͤ�9��9آ�9���9a��9���9���95��9w��9G��9��9@��9���9D��9��9���9
��9֢�9��9|��9���9���9���9��9��9͢�9x   x   ���9���9���9���9���9t��9���91��96��9��9
��9��9ƥ�9��9���9���9ƥ�9��9���9���9���95��9���9���9��9��9��9��9[��9��9x   x   s��9��9ã�9��99��9Ӧ�9[��92��9���9x��9���9��9���9Z��9;��9���9���9x��9���9���9���9��9i��9ģ�9���9��9���9*��9���9���9x   x   ١�9���9���9���9���9>��9���9��9}��9ߩ�9���98��9¨�9f��9%��92��9y��9У�9��9���9V��9-��9��9���9��9���9���9̤�9���9��9x   x   r��9���9l��9r��9Z��9M��9���9��9���9���9��9���9���9T��9���9r��9��9<��9@��9x��9��9&��9P��9q��9ަ�9&��9m��9��9���9���9x   x   t��9��90��9P��9i��9��96��9��9��99��9���9���9���9��9Ӥ�9ҟ�9���9���9ޤ�9Z��9"��9��9��9��9&��9$��96��9���9���97��9x   x   ���9 ��9"��9��9���9���9y��9ɥ�9��9���9��9���9���9���9��9���91��9��9\��9b��9���9���9���9���9���9_��9���9̤�9��9Ƥ�9x   x   ��9��9ר�9Ҥ�97��9��9H��9��9Z��9b��9T��9��9���9M��9��9��9���9o��9��9���94��9���9���9��9^��9��9���9���9ܥ�9Q��9x   x   ���9���98��9N��9��9ȥ�9��9���9<��9!��9���9դ�9��9ݤ�9��9���9H��9���9w��9ԣ�9��9 ��9���9���9*��94��9��9��9-��9��9x   x   ��9���9*��9���9���9p��9?��9���9���92��9r��9ӟ�9¦�9��9���9���9��9��9��9}��9���9���9Š�9i��9è�9>��9C��9��9���9��9x   x   p��9E��9!��9,��9u��9���9���9���9¦�9x��9��9���91��9Ħ�9I��9���9ȥ�9��9��9��9���9ͧ�9���9���9���9ʧ�9ѥ�9R��9��9��9x   x   ���9N��96��9l��9��9���9?��9��9��9ѣ�9=��9���9 ��9p��9���9��9��9��9��9~��9���9P��9���9���9���9��9���9'��96��9ߥ�9x   x   ���9��9��9���9c��9g��9��9���9���9��9>��9ݤ�9^��9��9y��9��9}��9��9@��9���9��9��9|��9Ǩ�9k��9L��9���9���96��9@��9x   x   ���9���9"��9���9���9��9���9��9���9���9y��9W��9d��9���9ӣ�9z��9��9~��9���9d��9���9Ϫ�9���9��9���9R��9s��9L��9m��9y��9x   x   X��9a��9&��9e��9d��9���9��9���9���9U��9��9!��9���93��9��9���9���9���9��9���9ݩ�9���9t��9��9���9���9	��9֤�9���96��9x   x   w��9��9���9V��9I��9��9բ�9:��9��9/��9&��9��9���9���9!��9���9Χ�9I��9��9̪�9���9/��9���9��9��9@��9E��9-��9Σ�9p��9x   x   i��9L��9!��9���99��9C��9��9���9g��9��9K��9���9���9���9���9Ƞ�9���9���9���9���9z��9Ȩ�9��9��92��9F��9Q��9���9M��9*��9x   x   Y��9���9 ��9$��9��9t��9{��9���9£�9���9p��9���9���9��9��9j��9���9���9ɨ�9��9	��9��9ߠ�9���9���95��9���9���9��9��9x   x   ���9��9���9���9ڥ�9���9���9��9���9��9��9(��9���9_��9)��9¨�9���9��9k��9���9���9��92��9���91��9���9z��9���9(��9��9x   x   b��9;��9���9%��91��9���9���9!��9��9���9&��9&��9Z��9��95��9<��9ʧ�9��9N��9O��9���9@��9E��9/��9���9���9e��9&��9���9���9x   x   i��9u��9��9'��9w��9���9���9��9���9���9m��98��9���9���9��9A��9̥�9���9���9t��9��9I��9Q��9���9y��9a��9%��9x��9͡�9��9x   x   ���9 ��9���9ʜ�9$��9n��9��9��9-��9Ф�9��9���9ͤ�9���9��9��9N��9#��9���9K��9Ӥ�9/��9���9���9���9'��9{��9k��9u��9ɢ�9x   x   H��9q��9-��9���9%��9���9��9\��9���9���9���9���9��9��9/��9���9��99��97��9p��9���9ѣ�9P��9��9'��9���9ˡ�9r��9~��90��9x   x   u��9��9O��9���9��9~��9Ң�9��9���9��9��95��9Ƥ�9S��9��9��9��9ߥ�9?��9x��93��9n��9)��9��9��9���9��9Ƣ�97��9ա�9x   x   ��9���95��9���9O��9���9���9 ��9���9���9���9���9���9���9��9���9���9j��9E��9��9���9��97��9l��9���9u��9���9"��9K��9���9x   x   ���9��9W��9���9���9i��9���9���9��9���9;��9)��9���9���9��9���9���9S��9���9J��9���9���9���9o��9���95��9:��9c��9,��9���9x   x   8��9V��9\��9���9d��9���9E��9���9���9���9���9��9j��9��9���9w��9��9��9.��9}��9���9���9���9>��9���9���9���9���9���9=��9x   x   ���9���9���9T��9%��9���9���9���9���92��9���9��9���9��9���9!��90��9Y��9���9���9��9���9?��9���9���9���9}��9���9|��9/��9x   x   O��9���9i��9'��9B��9���9���93��9���9&��9��9
��9���9_��9���9���9j��9_��9���9$��9���9a��9���9���9���9 ��9��9���9��9{��9x   x   ���9c��9���9���9���9���9p��9���9j��9���9���9e��9���9���9���9���9	��9���9��9v��91��9���9)��9:��9��9���9���9���9���9���9x   x   ���9���9D��9���9���9k��9��9���9���9���9���9Z��9���9���9���9���9
��9���9j��9���9���9���9���9���9���9���9���9%��9|��9���9x   x   ���9���9���9���93��9���9���9���9���9t��9��9U��9���9���9���9���9���9���9��9���9���9��9��9���9���9���99��9���9���9e��9x   x   ���9��9���9���9���9s��9���9���9���9��9���9I��9���9#��9���98��9���9���9���9z��9���9\��9���9���9G��9���9G��9���9s��9���9x   x   ���9���9���93��9!��9���9���9v��9��9���9���9-��9���9P��9���9f��9���9���91��9���9���9���9���9���9���9���9,��9���9��9���9x   x   ���9=��9���9���9��9���9���9��9���9���9���9!��9���98��9���9��9���9��9���9���9���9���9Z��9���9~��9���9L��9;��9���9y��9x   x   ���9*��9��9��9��9h��9Z��9T��9A��9-��9��9G��9d��9���9���9��9M��9���9z��9���9���9x��9���9���9���9��9"��9���9��9���9x   x   ���9���9m��9���9���9���9���9���9���9���9���9b��9���9���9��9���9���9+��9���9���9��9��9���9��9l��9G��9L��9���9���9���9x   x   ���9���9	��9��9a��9���9���9��9!��9S��9<��9���9���9���9!��98��9���9���9���9��9���93��9|��9���9��9~��9���9���9���9S��9x   x   ��9��9���9���9���9���9���9���9���9���9���9���9��9 ��97��9}��9���9t��9���9Z��97��9���9���9���9���9���9.��9���9-��9v��9x   x   ���9���9w��9#��9���9���9���9���99��9h��9��9��9���9;��9{��9f��9���9���9���9���9B��9���9��9���9Q��9y��9���9���9l��9���9x   x   ���9���9��91��9l��9	��9��9���9���9���9���9J��9���9���9���9���9��9���9���9v��9c��9���9���9l��9D��9���9���9���9���9;��9x   x   g��9W��9��9]��9Z��9���9���9���9���9���9��9���9+��9���9q��9���9���9���9w��9{��9���9���9���9���9T��9j��9���9X��9��9���9x   x   D��9���9.��9���9���9��9h��9��9���9,��9���9u��9���9���9���9���9���9z��9���9��9d��9���9���9���9���9\��9���9���9���9���9x   x   ��9N��9|��9���9&��9u��9���9���9{��9���9���9���9���9��9\��9���9x��9x��9��9��9��9���9O��9X��9��9���9���9:��9���9<��9x   x   ��9���9���9��9���9/��9���9���9���9���9���9���9��9���96��9B��9b��9���9f��9��9���9	��9
��9k��9���9���9���9��9	��9E��9x   x   ��9���9���9���9a��9���9���9!��9_��9��9���9w��9
��95��9���9���9���9���9���9���9��9��9��9���9���9���9���9���9]��9���9x   x   4��9���9���9>��9���9)��9���9��9���9���9`��9���9���9v��9���9��9���9���9���9N��9��9��9���9���9���9E��9���9&��9A��9���9x   x   m��9p��9=��9���9���9;��9���9���9���9���9���9���9��9���9���9���9n��9���9���9\��9j��9���9���9���9���9P��9��9���9���9��9x   x   ���9���9���9���9���9���9���9���9I��9���9{��9���9m��9#��9���9R��9C��9P��9���9��9���9���9���9���9���9��9v��9_��9��9���9x   x   v��97��9���9���9#��9���9���9���9���9���9���9��9E��9}��9���9y��9���9o��9Z��9���9���9���9F��9R��9#��9C��9��9���9)��9���9x   x   ���98��9���9~��9��9���9���98��9M��9*��9L��9%��9L��9���9-��9���9���9���9���9���9���9���9���9��9y��9��9B��9���9���9���9x   x   &��9b��9���9 ��9���9���9(��9���9���9���96��9���9���9���9���9���9���9[��9���9=��9��9���9$��9���9`��9���9���9���9���9���9x   x   O��9)��9���9y��9��9���9}��9���9u��9 ��9���9��9���9���9(��9m��9���9��9���9���9��9]��9?��9���9��9.��9���9���9���9���9x   x   ���9���9?��9,��9��9���9���9e��9���9���9{��9���9���9N��9r��9���91��9���9���99��9J��9���9���9��9���9���9���9���9���9o��9x   x   ��9��9�9$�9�9s�9K�9��9r�9.�9��9�9a�9&�9��9�9��9��9��9�9k�9��9��9�9-�9J�9��9��9k�9v�9x   x   ��9/	�9��9h�9t�9��9��9��9p�9-�9#�9��9-�9��9=�98�9H�9+�9�9��9�9��9a�9��9��9�9��9��9
�9{�9x   x   ��9��9��9*�9��9]�9��9��9��9��9��9�9��9e�9e�9��9��9�9[�9��9S�9��9T�9��9��9��9H�9��9��9m�9x   x   &�9j�9)�9�9�9��9S�9��9Y�9��9�9L�9��9"�9��9��9
�9��9�9��9��94�9�97�9G�9��9w�9p�9)�9i�9x   x   �9s�9��9�9e�9K�9�
�9J�9?�9��9�	�9��9�9��9��9��9	�9��9��9^�9��9#�9|�9��9O�9a�9��9��9��9�9x   x   q�9~�9`�9��9I�9}�9~�9��9��9��9��9t�9��9��9��9z�9\�9��9��9}�9!	�9��9��9��9	�9�9��9#�90�9,�9x   x   N�9��9��9W�9�
�9��9��9R�9�9X�9,�9��9��9P�99�9_�9��9��9��9��9��9��9G�9t�9��9��9t	�9��9�	�9��9x   x   ��9��9��9��9I�9��9M�9	�9��9#�97�9��9�9��9d�9l�9��9X�9�9!�9n�9��9��9��99�9��9r�9	�9;�9��9x   x   s�9o�9��9W�9<�9��9�9��9��9��9�9��9��9��9��9`�9P�9��9��9��9M�9��9H�9�9��9��93�9�9b�9�9x   x   2�9,�9��9��9��9��9U�9 �9��9H�9i�9��9��9��9��9�9��9v�9��9��9:�9��9�9�9L�9��9��9	�9��9�9x   x   ��9$�9��9�9�	�9��9,�9<�9�9i�9~�9��9�9z�9�9)�9�
�9�9��94�9Y�9��9��9��9��9e�9,�9U�9��9��9x   x   �9��9�9J�9��9v�9��9��9��9��9��9��9��9��9��9��9n�9\�9��9��9<�9<�9��9��9��9��9��9!�9e�9��9x   x   a�9-�9��9��9�9��9��9�9��9��9�9��9�94�9t�9��9q�9��9��9��9�9u�9��9��9��9��99�9y�9��9~�9x   x   $�9��9`�9 �9��9��9K�9��9��9��9x�9��97�9f�9�9��9��9��9x�9(�9�9��9[�9��9��9��9��9��9��9,�9x   x   ��9?�9d�9��9��9��96�9d�9��9��9 �9��9u�9�9�9��9��9��9��9�9�9��9��9-�9_�9U�9��9>�9U�9��9x   x   �9<�9��9��9��9~�9]�9k�9a�9
�9*�9��9��9��9��9��9��9�9N�9A�9��9��9��9��9��9��9<�9�9�9��9x   x   ��9E�9��9�9	�9]�9��9��9N�9��9�
�9k�9m�9��9��9��9v�99�9��9��9��9�9s�9��9��9��9��9;�9��9��9x   x   ��9-�9�9��9��9��9��9Y�9��9x�9�9a�9��9��9��9�99�9��9V�9��9��9��9��9�9P�9��9��9*�9��9`�9x   x   ��9	�9Z�9�9��9��9��9�9��9��9��9��9��9{�9��9K�9��9W�9Q�9�92�9��9�9��95�9W�9��9+�91�9��9x   x   �9��9��9��9]�9��9��9!�9��9��96�9��9��9)�9�9>�9��9��9�9��9��90�9��9�9��9��9�9+�9\�9��9x   x   j�9�9W�9��9��9	�9��9n�9L�98�9[�9=�9�9�9�9��9��9��9+�9��9��9��9~�9N�9��9W�9Y�9��9��9��9x   x   ��9��9��97�9 �9��9��9��9��9��9��9:�9s�9��9��9��9�9��9��97�9��9|�9��9�9��9��9��9}�9��9�
�9x   x   ��9`�9U�9�9��9��9G�9��9H�9�
�9��9��9�9]�9��9��9n�9��9�9��9|�9��9]�9��9��9F�9�9��9p�9��9x   x   �9��9��9:�9��9��9w�9��9�9�9��9��9��9��9,�9��9��9�9��9�9J�9�9�9��9S�98�9��9P�9%�98�9x   x   +�9��9��9F�9L�9�9��9=�9��9L�9��9��9��9��9[�9��9��9V�99�9��9��9��9��9S�9��9H�9��9�9��9��9x   x   G�9�9��9��9d�9�9��9��9��9��9f�9��9��9��9Y�9��9|�9��9V�9��9T�9��9B�94�9G�9��9�9`�9�9z�9x   x   ��9��9I�9s�9��9��9v	�9s�92�9��9-�9��9;�9��9��9;�9��9��9��9�9Y�9��9�9��9��9�9��9�9��9��9x   x   ��9��9��9n�9��9!�9��9
�9�9
�9U�9"�9|�9��9:�9�9:�9(�9*�9)�9��9~�9��9R�9�9c�9�9��9�9��9x   x   i�9
�9��9*�9��9-�9�	�9?�9b�9��9��9`�9��9��9W�9�9��9��9.�9W�9��9��9u�9'�9��9�9��9�9��9x�9x   x   s�9y�9m�9f�9�9(�9��9��9�9�9��9��9v�92�9��9��9��9b�9��9��9��9�
�9��9:�9��9y�9��9��9s�9��9x   x   �?�9C�9-A�9�?�9�D�9 A�9�B�9�B�9PB�9ZI�9�I�9�I�9 I�9KI�9�J�9cG�9J�97H�9hI�9cH�9�I�9�I�9JC�9QD�9�A�97@�9`D�9�@�9m@�9�B�9x   x   C�9�E�9�E�9�B�9qD�9�B�9?E�9I�9H�9�I�9F�9�H�9�F�9KK�9�F�9�F�9�L�9QF�9�H�9#G�9�I�9�G�9�F�9IE�9�C�9�D�9NB�9�F�9nF�99B�9x   x   .A�9F�9�F�9>�98H�9tH�9�E�9E�9�F�9
I�9�G�9�E�9�G�9xI�9�?�9�H�9�G�9�E�9G�9)H�9�F�9�F�9�F�9�G�9CG�9�>�9eF�9E�9	B�9�E�9x   x   �?�9�B�9>�9_>�9wG�9�B�9�D�9TE�97E�9(G�9�J�9NG�9�J�9MG�9H�9�J�9�G�9~J�9�G�9�F�9�C�9D�9�B�9jH�9 >�9�=�9�C�9�?�9�E�9�E�9x   x   �D�9uD�94H�9rG�9�@�9hF�9!J�9�G�9�G�9EI�9I�9�H�96J�9H�9(J�9�H�9�H�9�I�96F�9�G�9�K�9F�9�@�9�G�9VH�9_C�9�D�9=H�9lF�9iH�9x   x    A�9�B�9wH�9�B�9cF�9WI�9�D�9oB�9�E�9�E�9eF�9)H�9�F�9WF�9UH�9�F�9�E�9`F�9C�9�C�9wH�9�G�9�A�9�G�9�C�9�@�9�E�9�E�9�D�9�E�9x   x   �B�9;E�9�E�9 E�9 J�9�D�9�D�9�D�9H�9F�9;F�9*F�9�H�9�F�9�E�9�F�9BG�9�D�9�D�95E�9�I�9?D�9tG�9VD�9OB�9�H�9�C�9MD�9�D�9�H�9x   x   �B�9I�9E�9UE�9�G�9oB�9�D�9F�9�E�9�D�9�B�9\I�9�H�9 C�9WD�9#F�9TF�9�C�9�B�9�G�9�E�9�D�9�H�9iC�9uI�9mH�9�D�9�D�9�G�9:I�9x   x   PB�9 H�9�F�99E�9�G�9�E�9H�9�E�9{H�9nH�9�E�9�J�9�E�9�H�9H�9�E�9zH�9�F�9WF�9�D�9�G�9�G�9�B�9�C�9bC�9�D�9�G�9�D�96D�9�C�9x   x   XI�9�I�9	I�9)G�9GI�9�E�9F�9�D�9nH�9�H�9H�9�H�9'H�9�H�9�D�9�E�9fE�9RI�9nI�9^G�9�I�9J�9�I�9�F�9�E�9�D�9�D�9xE�9�E�9�J�9x   x   �I�9F�9�G�9�J�9I�9dF�99F�9�B�9�E�9H�9�E�9#H�9LF�9tB�9]F�95G�9LI�9"I�9"G�9�G�9�H�9>L�9LF�9
I�9�J�9+E�9�J�9HI�9$F�9�L�9x   x   �I�9�H�9�E�9LG�9�H�9(H�9&F�9UI�9�J�9�H�9$H�9�J�9�H�9�F�9�G�9�G�9�H�9�E�9�H�9�H�9�H�9GH�9�D�9{H�9�F�9
G�9gH�9�E�9fG�9H�9x   x   I�9�F�9�G�9�J�92J�9�F�9�H�9�H�9�E�9%H�9OF�9�H�9�H�9VF�9�K�9�I�9�F�9G�9�H�9.F�9cF�9�G�9F�9yE�9�H�9DE�98E�9�G�9�G�9+E�9x   x   NI�9HK�9}I�9SG�9H�9YF�9�F�9%C�9�H�9�H�9xB�9�F�9VF�9�G�9mG�9|J�9bK�9.I�92H�9�I�9�I�9�K�9yF�9�G�9�G�9�G�9�K�9�H�9.J�9'H�9x   x   �J�9�F�9�?�9H�9$J�9SH�9�E�9WD�9H�9�D�9_F�9�G�9�K�9iG�9L?�9bF�9�J�9I�9mF�9�I�9;I�9�K�9"I�9�H�9NH�9�J�9[J�9�H�9G�9�H�9x   x   bG�9�F�9�H�9�J�9�H�9�F�9�F�9$F�9�E�9�E�95G�9�G�9�I�9yJ�9_F�9�G�9K�9FG�9|G�9vJ�9rH�9SL�9�G�9>H�9KM�9�G�9�J�9�G�9�F�9�J�9x   x   !J�9�L�9�G�9�G�9�H�9�E�9CG�9RF�9|H�9dE�9KI�9�H�9�F�9cK�9�J�9K�9(J�9tJ�9^K�9�I�98I�9}M�9�J�9�L�9}I�9fI�9�K�9�I�9�J�9�K�9x   x   ;H�9QF�9�E�9J�9�I�9aF�9�D�9�C�9�F�9QI�9!I�9�E�9 G�9.I�9I�9HG�9zJ�9�H�9BH�9�E�9�D�9M�9�M�9�C�9FF�9kH�9I�9�J�9�E�9�I�9x   x   gI�9�H�9G�9�G�95F�9C�9�D�9�B�9UF�9pI�9G�9�H�9�H�9.H�9iF�9}G�9cK�9DH�9�N�9�J�9]H�9VK�9�H�9�J�9]N�9�G�9K�9�G�9�F�9�H�9x   x   dH�9G�9*H�9�F�9�G�9�C�93E�9�G�9�D�9`G�9�G�9�H�9,F�9 J�9�I�9wJ�9�I�9�E�9�J�9J�9G�9nF�9^J�9�J�9�F�9�J�9�I�9OJ�9�H�9�E�9x   x   �I�9�I�9�F�9�C�9�K�9yH�9�I�9�E�9�G�9�I�9�H�9�H�9gF�9�I�9>I�9sH�9:I�9D�9_H�9G�9DE�9�F�9`H�9QD�9�G�9KI�9�H�9_J�9�G�9�H�9x   x   �I�9�G�9�F�9D�9F�9�G�9<D�9�D�9�G�9J�9<L�9KH�9�G�9�K�9�K�9OL�9�M�9M�9[K�9eF�9�F�9NK�9LM�9wN�9�L�9�K�9QK�9G�9|G�9�K�9x   x   LC�9�F�9�F�9�B�9�@�9�A�9sG�9�H�9�B�9�I�9NF�9�D�9F�9{F�9#I�9�G�9�J�9�M�9�H�9\J�9dH�9RM�9hI�92H�9H�9TG�9�F�9�D�9wG�9�I�9x   x   LD�9GE�9�G�9gH�9�G�9�G�9ZD�9fC�9�C�9�F�9	I�9wH�9uE�9�G�9�H�9AH�9�L�9�C�9�J�9|J�9PD�9wN�9.H�9�H�9AH�9�C�9�H�9xH�9 F�9MC�9x   x   �A�9�C�9CG�9&>�9[H�9�C�9QB�9tI�9_C�9�E�9�J�9�F�9�H�9�G�9KH�9KM�9�I�9GF�9ZN�9�F�9�G�9�L�9H�9GH�9{I�9[G�9�J�9�E�9vD�9�H�9x   x   7@�9�D�9�>�9�=�9bC�9�@�9�H�9mH�9�D�9�D�9+E�9G�9BE�9�G�9�J�9�G�9fI�9kH�9�G�9�J�9KI�9�K�9SG�9�C�9\G�90D�9ME�9�C�9�H�9lI�9x   x   ^D�9TB�9cF�9�C�9�D�9�E�9�C�9�D�9�G�9�D�9�J�9fH�94E�9�K�9[J�9�J�9�K�9!I�9K�9�I�9�H�9OK�9�F�9�H�9�J�9ME�9�G�9�D�9C�9�F�9x   x   �@�9�F�9E�9�?�9=H�9�E�9LD�9�D�9�D�9yE�9GI�9�E�9�G�9�H�9�H�9�G�9�I�9�J�9�G�9PJ�9_J�9G�9�D�9{H�9�E�9�C�9�D�94E�9E�9�G�9x   x   m@�9qF�9B�9�E�9nF�9�D�9�D�9�G�9/D�9�E�9!F�9fG�9�G�92J�9G�9�F�9�J�9�E�9�F�9�H�9�G�9yG�9pG�9�E�9sD�9�H�9C�9E�9�F�9�E�9x   x   �B�98B�9�E�9�E�9kH�9�E�9�H�9:I�9�C�9�J�9�L�9H�9+E�9(H�9�H�9�J�9�K�9�I�9�H�9�E�9�H�9�K�9�I�9OC�9�H�9iI�9�F�9�G�9�E�9rF�9x   x   �{�9|�9�{�9}}�9^}�9�~�9��9���9��9w|�9h~�9�~�9���9���9��9��9��9H��9���9k~�9~�9�|�9��9���9��9�~�9�}�9<~�9Hz�9�{�9x   x   |�9�}�9]z�9k}�9��9��9x��9}�9�}�9{�9�9
��9���9/~�9��9҂�9�~�9n��9;��9�~�9n{�9^~�9�|�9���9��9@�9�|�9T{�9�~�9�{�9x   x   �{�9]z�9#{�9H��9\z�9�z�9�|�9��9���9L�9Z��9��9n��9��9҄�9���9>��9��9���9m�9��9��9�|�9�y�9�z�9��9Jz�9�y�9z{�9{�9x   x   {}�9g}�9I��9��9~~�9�~�9N�9�}�9���9�{�9~�9^~�9�}�9��9���9�}�9�~�9�}�9�{�9���9~�92�9I�9�~�9��9ۂ�9~�9�}�9m�9�~�9x   x   ^}�9��9`z�9�~�9Ӂ�9�~�9E}�95��9U��95|�9��9��9~�9���9�}�9��9ׄ�9X|�9Ā�9t��9�|�9�~�9v��97�9�z�9�~�9}�9cz�9�v�9_{�9x   x   �~�9��9�z�9�~�9�~�9�|�9�~�9@��9��9g}�9���9}�9Y��91��9�}�9r��9�}�9h��9��9�~�9l}�9m�9o~�9kz�9��9L�9�|�9�y�9Cy�9
|�9x   x   ��9u��9�|�9O�9F}�9�~�9d��9���9/�9]�9���9��9���9&��9#��9Z�93~�9���9~��9�~�9B|�9r�9-}�9Z��9��9�{�9Հ�9ށ�9#��9�|�9x   x   ���9}�9��9�}�94��9?��9���9��9��9o��9���9��9��9���9���9Ã�9��9t��91��9���9z~�9f�9}�9���9{y�9J}�9�|�9z}�9�|�9�x�9x   x   ��9�}�9���9���9U��9��90�9��9+��9�~�9ހ�9�}�9*��9�~�9��9N��9�~�9/��9��9Ԁ�9X��9�}�9��9���9k|�9��9�|�9���9�|�9��9x   x   v|�9{�9L�9�{�95|�9f}�9_�9n��9�~�9�~�9��9��9�~�9m�9���9=�9s}�9Q|�9c|�9�9�{�9�|�9���9D��9"��9K��9!��9��9Ł�9t��9x   x   k~�9�9X��9~�9��9���9��9���9ހ�9��9[��9��9#��9���9%��9ʃ�9��9}}�9P��9~�9�}�9E|�9,{�94~�9�~�9��9�~�9}�9�{�9 }�9x   x   �~�9��9��9`~�9%��9}�9��9��9�}�9��9��9�~�9��9��9L}�9��9"�9b��9���9�~�9���9}��9���9܀�9���9���9n��9)��9���9�~�9x   x   ���9���9l��9�}�9~�9S��9���9��9&��9�~�9 ��9��9���97��9~�9�}�9��9܁�9(��9��9E�9���9��9ʄ�9���91��9Q��9���9���9���9x   x   ���90~�9��9��9���9'��9*��9��9�~�9l�9���9��96��9L��9���9g��9;~�9(��9���9Ȃ�9���9�~�9��9��9���9���9��9}��9��9 ��9x   x   ��9��9̈́�9���9�}�9�}�9"��9���9��9���9)��9I}�9~�9���9���9Q��9G��9��9`��9u��9��9}��9���9y��9݅�9Q��98��9e��9��9Q��9x   x    ��9ӂ�9���9�}�9��9p��9[�9�9N��9<�9̓�9��9}�9i��9O��9P��9L��9V��9��9��9q~�9���9���9���9��9f~�9Ё�9g��9g��9��9x   x   
��9�~�9@��9�~�9ڄ�9�}�95~�9
��9�9s}�9��9 �9��9>~�9L��9Q��9Ɓ�9J��9���97��9
��9)��9p�9N��9z��9u��9X��9=��9 ��9��9x   x   E��9k��9��9�}�9V|�9d��9���9p��9(��9Q|�9~}�9a��9ځ�9#��9��9V��9B��9[��9Յ�9��9O��9
��9��9~��9U��9��9���9ق�9���9	��9x   x   ���9:��9���9�{�9���9��9���94��9��9h|�9Q��9���9-��9���9`��9��9���9Ӆ�9���9҂�9��9��9L��9#��9<��9��9͂�9���9X��9X��9x   x   j~�9�~�9p�9���9x��9�~�9�~�9���9Ԁ�9�9~�9�~�9��9̂�9u��9��97��9
��9ւ�9���9���9���9��9���9���9���9w��9��9���9���9x   x   ~�9q{�9��9~�9�|�9i}�9@|�9|~�9U��9�{�9�}�9���9@�9���9���9o~�9��9K��9 ��9���9���9���9���9^��9ޅ�9|~�9���9t��9��9��9x   x   �|�9[~�9��90�9�~�9k�9q�9j�9�}�9�|�9B|�9~��9���9�~�9���9���91��9
��9��9���9���9\��9r��9���9V��9K��9�9���9ځ�9�|�9x   x   ��9�|�9�|�9O�9x��9q~�91}�9}�9��9���9){�9 ��9��9��9���9���9q�9��9N��9��9���9m��9��9���9Å�9e��9׃�9���9�|�9���9x   x   ���9���9�y�9�~�97�9nz�9Y��9���9���9C��93~�9߀�9Ʉ�9��9y��9���9R��9{��9'��9���9^��9���9���9���9~��9.��9��9�|�9���9���9x   x   ��9��9�z�9��9�z�9��9��9{y�9j|�9"��9�~�9���9��9���9݅�9��9|��9T��9?��9���9ޅ�9T��9Ņ�9{��9���9��9_�9́�9x|�9nx�9x   x   �~�9:�9��9ۂ�9�~�9M�9�{�9G}�9��9O��9��9���9-��9���9Q��9c~�9v��9��9��9���9}~�9I��9f��9,��9��9x~�9���9Á�9	}�9�|�9x   x   �}�9�|�9Lz�9~�9}�9�|�9ր�9�|�9�|�9 ��9�~�9s��9R��9��98��9с�9S��9���9˂�9w��9���9�9ڃ�9��9_�9���9�{�9�}�9r��9o|�9x   x   =~�9Q{�9�y�9�}�9`z�9�y�9��9y}�9���9��9}�9,��9���9y��9h��9e��99��9܂�9���9��9r��9���9��9�|�9΁�9�9�}�9���9�y�9Hz�9x   x   Jz�9�~�9z{�9j�9�v�9Gy�9#��9�|�9�|�9ȁ�9�{�9���9���9��9��9h��9��9���9W��9���9��9ށ�9�|�9���9~|�9}�9p��9�y�9w�9�~�9x   x   �{�9�{�9#{�9�~�9[{�9|�9�|�9�x�9��9p��9}�9�~�9���9��9Q��9��9��9	��9S��9���9��9�|�9���9���9mx�9�|�9l|�9Hz�9�~�9�|�9x   x   ���93��9=��9O��9���9���9���9��9���9���9Z��9���9���9���9���9��9���96��9w��9	��9���9��9��9{��9l��9��9g��9Ҹ�9��9��9x   x   3��9[��9>��9ɵ�9z��9��9���9@��9H��9'��9��9׶�9���9���9L��9���9��9y��9��9i��9{��9c��9��9ٶ�9���9���9���9��9���9���9x   x   ;��9>��9x��9ҵ�9H��9��9l��9��9?��9��9���9Ƽ�9��9[��9���9չ�9;��9x��9���9���9���95��9��9��9ĳ�9m��9��9���9/��9��9x   x   N��9˵�9ӵ�9��9���9f��9���9R��9���9��9��9_��9��9Y��9���9���9q��9���9Ž�9���9׹�9C��94��9���9+��9���9���9h��9��9���9x   x   ���9x��9H��9���9!��9���96��9Ƕ�9��9���9��9��9��91��9���9��9���9��9��9���9h��9���9A��9`��9	��9��9D��9��9���9��9x   x   ���9��9��9a��9���9���9���9R��9e��9���92��9���9λ�9��9��9��9ɼ�9��9˵�9_��9���9���9���9��9��9���9��9���9��9ƶ�9x   x   ���9���9l��9~��98��9���9]��9·�9Ȼ�9��9K��9 ��9��9۹�9��9p��9���9ٷ�9��9Y��9>��90��9V��9���9¶�9��9���9��9���91��9x   x   ��9>��9��9P��9˶�9Q��9÷�9G��9���9���9z��9ָ�9��9g��9���9���9J��9���9��9B��9���9��9��9��9���97��9���9���9A��9b��9x   x   ���9G��9?��9���9��9]��9Ļ�9���9���9T��98��9 ��9Q��9���91��9N��9ĺ�9A��9Y��9���9`��9���9���9D��9���9���9���9;��9ȹ�9p��9x   x   ���9'��9��9��9���9 ��9	��9���9V��9���9���9���9���9ͻ�9���9Ż�9q��9���9B��9Ⱥ�9Ż�9���9���9���9:��9��9.��9]��9z��9A��9x   x   V��9��9���9��9��90��9M��9w��9:��9���9���9}��9��9���9���9Ʒ�9k��9���9��9=��9���9ƹ�9
��9��9���9���9���9N��9���9M��9x   x   ���9ٶ�9ȼ�9`��9��9���9��9ϸ�9#��9��9y��9̻�9(��9��9"��9���9��9���9���9���9���9��9'��9��9\��9���9`��9���9A��92��9x   x   ���9���9��9��9��9ͻ�9��9��9T��9���9��9,��91��9I��9��9��9&��9���9���9Ƚ�9���9���9=��9���9͹�9 ��9���9���9d��9���9x   x   ���9���9_��9X��95��9���9ܹ�9h��9���9ͻ�9��9��9M��9 ��9"��9J��9|��9���9Ⱥ�9��9���9~��97��9��9���9��9P��9;��9��9��9x   x   ���9M��9���9���9���9��9��9���91��9���9���9%��9��9"��9½�9���9���9,��9˼�9(��9E��9��9���9���9���9��9��9���9��9��9x   x   ��9���9չ�9���9��9��9s��9���9L��9���9ķ�9���9��9G��9���9D��9��9z��9���9 ��9Q��9%��9G��9���9O��9���9$��9���9��9���9x   x   ���9��9=��9r��9���9˼�9���9G��9Ⱥ�9r��9j��9��9&��9~��9���9��9#��9Ƽ�9���9��9���9���9P��9׺�9���9���9��9[��9���9��9x   x   7��9z��9y��9���9��9��9׷�9���9F��9���9~��9���9���9���9)��9z��9ü�9���9���9���9���9,��9���9��90��9l��9]��9��9]��9���9x   x   w��9��9���9Ž�9��9ȵ�9��9��9[��9>��9��9���9���9ʺ�9̼�9���9 ��9���9i��9��9ɾ�9^��9���9t��9U��9U��9ݽ�9��9���9��9x   x   ��9d��9���9���9���9b��9Y��9>��9���9ú�9:��9���9ƽ�9��9&��9���9��9���9��9���9���9���9:��9о�9U��9���9���9��9A��9ƾ�9x   x   ���9|��9���9ӹ�9k��9���9=��9���9`��9ƻ�9���9���9���9���9D��9Q��9���9���9ľ�9���9K��9���9���9Q��9��9���9���9��9Ҽ�9%��9x   x   ��9g��95��9@��9���9���91��9��9���9���9ʹ�9��9���9~��9��9&��9���91��9^��9���9���9���9��9ݹ�9��9���9���9���9/��9���9x   x   ��9��9���97��9B��9���9P��9��9���9���9
��9"��9=��93��9���9G��9P��9���9���92��9���9߽�9r��9��9���9W��9Ϻ�9P��9���9��9x   x   {��9ض�9��9}��9_��9��9|��9���9>��9���9��9��9���9��9���9���9ֺ�9��9r��9ξ�9W��9߹�9��9���9V��9��9{��9���91��9˸�9x   x   k��9���9Ƴ�9(��9	��9��9���9���9���9:��9���9Y��9̹�9���9���9M��9���90��9T��9P��9��9��9���9Q��9
��9���9R��9���9���9`��9x   x   ��9���9q��9���9��9���9��9<��9���9��9���9���9��9��9��9���9���9l��9T��9���9���9���9X��9��9���9���9���9���9=��9���9x   x   j��9��9��9���9A��9#��9���9���9���9.��9���9a��9���9R��9��9"��9"��9^��9ݽ�9���9ÿ�9���9Һ�9w��9Q��9���9��9���90��9>��9x   x   Ҹ�9��9���9i��9��9���9��9���97��9[��9L��9���9���9?��9���9���9Z��9	��9��9��9��9���9P��9���9���9���9���9��9w��9M��9x   x   ��9���91��9��9���9޺�9���9C��9ȹ�9}��9���9@��9d��9��9��9��9���9_��9���9C��9Ѽ�9.��9���93��9��99��9/��9x��9���9���9x   x   ��9���9��9���9��9ȶ�94��9e��9m��9=��9Q��93��9���9��9��9���9��9���9��9Ⱦ�9!��9���9��9˸�9`��9���9=��9O��9���9[��9x   x   X��9���9G��9���9a��9���9���95��9���9E��9��9���9���9���9���9���9���9���9F��9���9���9���9^��9���9���9���9���9���9���9���9x   x   ���9��9���9���9���9���9��9���9^��9]��9���9W��9���9���9c��9���9���9���9���9���9���9���97��9���9��9��93��9���9���9m��9x   x   F��9���9I��9��9V��9���9��9B��9���9��9v��9]��9���9���9���9���9���9'��9B��9���9f��9���9��9/��9>��95��9}��9���9��9n��9x   x   ���9���9��9���9���9���9���9���9?��9���9B��9��9��9���9��95��9S��9���9���9���9���9���97��9���9���9u��9���9U��9���9.��9x   x   _��9���9U��9���9���9���9���9���9���9���9���9���9���9���93��9a��9P��9e��9���9a��9���9v��9���9 ��9���9��9B��9���9���9���9x   x   ���9���9���9���9���9���9���9N��9���9���9K��9��9���9N��9d��94��9���9i��9��9��9p��9���9���9���9���9M��9���9Q��9���9���9x   x   ���9��9��9���9���9���9X��9b��9���9���9Y��9K��9���9���9���9���9���9T��9���9��9?��9[��9���9���9���9���9���9b��9���9���9x   x   4��9���9E��9���9���9N��9i��9-��9���9���9���9&��9���9���9���9%��9���9���9��9G��9���9���9F��9���9���9���9��9���99��9&��9x   x   ���9_��9���9>��9���9���9���9���9��9z��9���9w��9L��9$��9��9T��9���9+��9���9M��9��9t��9���9v��9���9��9���9?��9��9���9x   x   G��9]��9��9���9���9���9���9���9x��9"��9��9��9���9x��9���9���9@��9���9b��9��9���9{��9��9���9���9��9p��9���9���9u��9x   x   ��9���9u��9=��9���9N��9[��9���9���9��9���9���9��9���9f��98��9'��9k��9���9���9���9y��9��9X��9��9E��9���9k��9���9s��9x   x   ���9R��9[��9��9���9��9K��9%��9z��9��9���9���9���9���9:��98��9���9���9���9A��9l��9'��9��9|��9��9���9���9
��9���9;��9x   x   ���9���9���9��9���9 ��9���9���9M��9���9��9���9c��9���92��9&��9	��9���9��9U��9���9���9���9���9���9_��9i��9|��9U��9���9x   x   ���9���9���9���9���9Q��9���9���9��9v��9���9���9���9���9+��9:��9���92��9���9'��9Q��9���9���9���9��9���9��9���9���9���9x   x   ���9]��9���9��9.��9b��9���9���9 ��9���9c��97��9+��9+��9w��9���9G��9���9X��9d��9���9���9'��9���9
��9���9���9F��9���9u��9x   x   ���9���9���9;��9b��97��9���9*��9V��9���97��9=��9(��9<��9���9��9n��9���9���9���9g��9(��9'��9��9���9���9���9��9Q��9���9x   x   ���9���9���9X��9L��9���9���9���9���9@��9#��9���9��9���9H��9n��9o��9���9\��9E��9l��9I��9��9���9���9��91��9��9���9���9x   x   ���9���9$��9���9c��9j��9X��9���9)��9���9m��9���9���97��9���9���9���9��9#��9���9���9���9���9���9h��9���9���9���9b��9���9x   x   E��9���9A��9���9���9��9���9��9���9c��9���9���9��9���9T��9���9\��9!��9���9���9���9���9���9  �9��9F��9P��9���9���9���9x   x   ���9���9���9���9_��9��9{��9F��9Q��9��9���9F��9V��9'��9c��9���9A��9���9���9���9��9��9���9���9���9��9���9���9B��9���9x   x   ���9���9h��9���9���9p��9B��9���9��9���9���9n��9���9R��9���9j��9l��9���9���9���9���9���9���9h��9?��9.��9���9��9��9���9x   x   ���9���9���9���9u��9���9`��9���9r��9v��9s��9%��9���9���9���9'��9D��9���9���9��9���9���9w��9A��9���9���9���9=��9L��9e��9x   x   ]��9:��9��99��9���9���9���9I��9���9��9��9��9���9���9&��9.��9��9���9���9���9���9t��9��9���9D��9c��9���9���9���9I��9x   x   ���9���9/��9���9#��9���9���9���9q��9���9X��9x��9���9���9���9��9���9���9 �9���9l��9A��9���9���9���9���9���9���9���9���9x   x   ���9��9B��9���9���9���9���9���9���9���9��9��9���9��9	��9���9���9e��9��9���9>��9���9D��9���9��9���9e��9{��9���9%��9x   x   ���9��91��9s��9��9I��9���9���9��9��9F��9���9f��9���9���9���9��9���9H��9��90��9���9f��9���9���9���9���9��9~��9���9x   x   ���97��9y��9���9C��9���9���9��9���9s��9���9���9i��9���9���9���97��9���9R��9���9���9���9���9���9f��9���9 ��9n��9���9���9x   x   ���9���9���9T��9���9O��9f��9���9A��9���9l��9��9��9���9H��9��9��9���9���9���9��9>��9���9���9{��9��9o��9���9��9p��9x   x   ���9���9���9���9���9���9���96��9��9���9���9���9W��9���9���9O��9���9[��9���9?��9��9L��9���9���9���9��9���9��9���9���9x   x   ���9q��9l��9,��9���9���9���9&��9���9z��9p��9;��9���9���9p��9���9���9���9���9���9���9g��9F��9���9&��9���9���9r��9���9���9x   x   �/�9�,�9x)�9_,�9W-�9�,�9�1�9#1�9)0�990�9�3�9�3�95�9X2�9�0�9�4�9�2�9�3�94�9�4�9U2�9#1�9V0�9�.�9�2�9�-�9�,�9�+�9}+�9-�9x   x   �,�90�9�(�9H+�9/-�9�,�90�9�0�9m/�9�5�9�4�96�902�95�96�9n5�9�2�9?2�9^6�9"5�9�5�92.�93�9�/�9�+�9�-�9�+�9$(�9o.�9�,�9x   x   y)�9�(�9�,�9I.�9U*�9-)�91�9�1�9�5�9�5�9�4�9�6�93�9�6�9+3�9�8�9�4�9�6�9�3�96�9q6�9R0�9�0�9*�9*�9�-�92-�9<)�9�*�9�&�9x   x   [,�9F+�9I.�9+�9�,�9G.�9'2�9r/�9�1�9=1�9�2�96�9�3�995�9�3�9�2�9�4�9U4�92�9l/�9k1�9�2�9�-�9�,�9�+�9/.�9�*�9�+�9B,�9�-�9x   x   W-�91-�9U*�9�,�9�1�90�9�.�9�/�9�2�9�1�94�9�1�960�9a;�9a1�9�3�964�9�/�9j4�9&/�95-�9�0�9�1�9�,�9�)�9�-�9�-�9�.�9�(�9�-�9x   x   �,�9�,�9-)�9G.�90�9�,�9 0�9�5�9�2�9$2�9Q5�9�1�9�3�9[4�9�/�9�4�9}3�9�1�9�5�91�9Q-�9�/�9�.�94)�9P,�9,�9{+�9c,�9,�9,�9x   x   �1�90�91�9&2�9�.�90�9/1�91�9�0�9�0�9e2�94�9�2�9�3�9_4�9|/�9�1�91�9�0�9�/�9�.�9<2�90�9 1�92�9�-�9#0�9=2�9�0�9�,�9x   x   (1�9�0�9�1�9u/�9�/�9�5�91�9�2�9�1�9�4�9p5�9A0�9~0�9
5�9�4�91�9<2�9�1�96�9�/�9Y/�9�2�9�0�9	0�9,�9�,�9�,�9',�9�,�9�,�9x   x   +0�9j/�9�5�9�1�9�2�9�2�9�0�9�1�9�-�9Q3�95�9Z2�9�5�9�1�9J/�9D2�9+0�92�9�2�9�1�9�4�95/�9�0�9�2�9�1�9�.�9-�9!/�9e2�9C1�9x   x   70�9�5�9�5�9;1�9�1�9#2�9�0�9�4�9O3�985�9�4�9]3�97�9�3�9#2�9d1�9�2�9�1�9>0�9�6�9�5�9L0�9�2�983�9f5�9>3�9�3�9�3�9�3�94�9x   x   �3�9�4�9�4�9�2�94�9V5�9e2�9s5�95�9�4�9�3�9�4�9E3�9�6�94�9�3�9�3�9l4�9�4�9�3�9�3�9�2�9&.�9D-�9[/�9l+�90�9�-�9h-�9�2�9x   x   �3�96�9�6�9 6�9�1�9�1�94�9F0�9Z2�9a3�9�4�9�2�9�0�9�2�91�9#4�9m4�9q6�9�6�9L4�9u8�9o7�9+7�9�7�9�5�9�4�9�7�97�9v7�9B9�9x   x   5�942�93�9�3�950�9�3�9�2�90�9�5�97�9A3�9�0�9q2�9�4�9B/�9u3�9x4�992�994�9M4�9U5�9d4�9o7�9J3�9I6�9�3�9�6�9�5�9�4�9A4�9x   x   V2�9#5�9�6�945�9`;�9Z4�9�3�95�9�1�9�3�9�6�9�2�9�4�9�;�9�4�9�6�9�3�9�2�9�8�9�3�9"2�9O6�96�9;4�9v4�9D6�9�5�9�1�94�9(8�9x   x   �0�96�9,3�9�3�9c1�9�/�9]4�9�4�9L/�9!2�94�91�9E/�9�4�9[3�9�5�922�9z7�9�;�9�7�9�7�9[7�9�9�9H8�9�8�98�9�7�9b8�9�;�9�7�9x   x   �4�9q5�9�8�9�2�9�3�9�4�9z/�91�9A2�9g1�9�3�9!4�9s3�9�6�9�5�9�4�95�9Q5�997�9[9�9�5�9�8�9:6�9c7�9b8�9%5�9m9�9
6�9�5�9`6�9x   x   �2�9�2�9�4�9�4�944�9}3�9�1�9<2�9*0�9�2�9�3�9i4�9x4�9�3�902�95�9p;�9�7�98�9�9�9D:�9`:�9�3�9�:�9�:�9>:�9�8�9%9�9X9�9�4�9x   x   �3�9E2�9�6�9\4�9�/�9�1�9	1�9�1�92�9�1�9n4�9n6�9?2�9�2�9{7�9P5�9�7�9�3�9F9�9�;�9�:�9�:�9r9�9�:�9;�9�8�9�2�98�9�7�9|6�9x   x    4�9[6�9�3�92�9i4�9�5�9�0�96�9�2�9@0�9�4�9�6�994�9�8�9�;�967�98�9G9�9�7�9j3�98�94�919�9?3�9�8�9�:�98�9�5�9�:�9r8�9x   x   �4�9!5�96�9j/�9,/�91�9�/�9�/�9�1�9�6�9�3�9L4�9M4�9�3�9�7�9\9�9�9�9�;�9i3�9=�9s:�9T:�9<�9x3�9�9�9_9�9�:�9�7�95�9�3�9x   x   [2�9�5�9n6�9i1�93-�9R-�9�.�9T/�9�4�9�5�9�3�9t8�9R5�92�9�7�9�5�9G:�9�:�98�9s:�9	<�9t:�9�8�9�;�9<�94�9�7�9G1�9D4�9f9�9x   x   &1�90.�9N0�9�2�9�0�9�/�9;2�9�2�95/�9P0�9�2�9r7�9c4�9M6�9Z7�9�8�9e:�9�:�94�9U:�9p:�9R4�9\9�9�8�9k9�9<8�9�6�9U5�9�7�9	3�9x   x   Y0�93�90�9�-�9�1�9�.�90�9�0�9�0�9�2�9#.�937�9n7�9%6�9�9�986�9�3�9m9�919�9&<�9�8�9X9�9�6�96�9�9�9?5�97�9�6�9 -�9M3�9x   x   �.�9�/�9*�9�,�9�,�94)�91�90�9�2�923�9F-�9�7�9D3�9?4�9E8�9a7�9�:�9�:�9:3�9s3�9�;�9�8�96�9�8�9j4�9|4�9Q7�9�.�9�3�9G2�9x   x   �2�9�+�9!*�9�+�9�)�9M,�92�9�,�9�1�9f5�9\/�9�5�9E6�9v4�9�8�9a8�9�:�9;�9�8�9�9�9<�9m9�9�9�9h4�9�5�95�9�.�9 4�91�9	/�9x   x   �-�9�-�9�-�9/.�9�-�9,�9�-�9�,�9�.�9<3�9h+�9�4�9�3�9G6�9�8�9$5�9@:�9�8�9�:�9b9�94�9>8�9<5�9w4�95�9�,�983�9�0�9F+�9>+�9x   x   �,�9�+�94-�9�*�9�-�9|+�9%0�9�,�9
-�9�3�90�9�7�9�6�9�5�9�7�9i9�9�8�9�2�98�9�:�9�7�9�6�97�9O7�9�.�953�9�+�9m,�93�9Z+�9x   x   �+�9#(�9:)�9�+�9�.�9f,�9<2�9!,�9"/�9�3�9�-�97�9�5�9�1�9k8�96�9%9�9!8�9�5�9�7�9I1�9V5�9�6�9�.�94�9�0�9f,�9�0�9�+�9�.�9x   x   ~+�9l.�9�*�9E,�9�(�9,�9�0�9�,�9k2�9�3�9e-�9x7�9�4�9 4�9�;�9�5�9Y9�9�7�9�:�95�9D4�9�7�9�,�9�3�91�9L+�93�9�+�9�(�9�,�9x   x   -�9�,�9�&�9�-�9�-�9,�9�,�9�,�9E1�94�9�2�9E9�9C4�9+8�9�7�9c6�9�4�9�6�9u8�9�3�9j9�93�9P3�9B2�9/�9:+�9Y+�9�.�9�,�9�%�9x   x   �g�9Dd�9�g�9�j�9
j�9k�9mo�9<k�9!p�9q�9�t�97p�94r�9�v�92u�9by�9�v�9]w�9[q�9 q�9,t�9Ur�9�o�9Yi�9�o�9�k�9�i�9j�9k�9�d�9x   x   Hd�9�i�9�i�9Gg�9h�9�l�9�i�9�j�9�p�94o�9n�9@n�9�t�9�u�9�s�9�r�9�s�9�u�9�m�90n�9�n�9}o�9�l�9�i�9�l�9�g�9dh�9�h�9�f�9d�9x   x   �g�9�i�9�h�9�i�9�m�9�n�9�m�9]l�9�k�9�k�96p�9Or�9�r�9ur�9*p�9t�9_s�9Rr�9�o�9�k�9�l�9kk�91m�9�o�9/m�9�h�9>i�9{j�9j�9f�9x   x   �j�9Ig�9�i�9�l�9'm�9To�9�n�9�n�9np�9}t�9to�9q�9Lu�9�q�9gp�9�t�9{o�9sp�9�t�9o�9�o�9�n�9o�9Gl�9Mn�9Si�9�f�9#j�9�g�9Uj�9x   x   
j�9h�9�m�9%m�9�i�9j�9Pp�9Am�95o�99r�9 o�9�s�9�r�9�o�9s�9�u�9|o�9Xp�9�p�9�l�9�o�9mj�9�j�9�l�9�l�9Xi�9Cj�9fj�9�h�9)i�9x   x   k�9�l�9�n�9Qo�9j�9Ds�9As�9m�9Zq�9�s�9 r�9hv�9�r�9�s�9Yt�9�p�9u�9q�96l�9�s�9Ws�9�h�9"p�9o�9nl�9�i�94h�9�n�9�m�9�h�9x   x   po�9�i�9�m�9�n�9Pp�9Hs�9�m�98n�9it�9#q�9^m�9kr�9;r�9qr�9�o�9p�9�t�9pn�9�m�9�r�9�q�9Bn�9�l�9k�9Go�9�k�9�i�97f�9Tk�9-j�9x   x   9k�9�j�9_l�9�n�9;m�9 m�95n�9q�9It�98t�9+q�9Zs�9�r�9)p�9 t�9+t�9�p�9jn�9%m�9�l�9n�9�m�9j�9j�9�k�9:s�9Fn�9�l�9�r�9�k�9x   x   p�9�p�9�k�9np�97o�9[q�9gt�9Lt�9p�9�p�9or�9*s�9It�9�o�9Fq�9�t�9;t�9�p�9cp�9�p�97k�9ep�9q�9Ym�9Ql�9<o�9�n�9to�9n�9�k�9x   x   q�96o�9�k�9zt�98r�9�s�9'q�99t�9�p�9zq�9�p�9�n�9]r�9�q�9�q�97q�9�t�9zq�9Ys�9�l�9�n�96q�9�m�9�p�9�n�9�o�9Vq�9�l�9Op�9�o�9x   x   �t�9n�95p�9to�9�n�9 r�9_m�9)q�9mr�9�p�94q�9_p�9q�9:r�9�o�9;p�9�n�9q�9�o�9�m�9ou�9n�9t�9�r�9�q�9�u�9r�9�s�9�s�9�m�9x   x   8p�9>n�9Ir�9q�9�s�9fv�9lr�9Us�9(s�9�n�9\p�9t�9#s�9wp�9�u�9�u�9�o�9�q�9un�9p�9�p�9ep�9Fv�9vo�9uu�9�s�9�o�9�u�9�o�95r�9x   x   4r�9�t�9�r�9Mu�9�r�9�r�9<r�9�r�9Ht�9\r�9 q�9's�9�s�9Ns�93r�9�t�9zs�9fu�9r�9Qt�9�u�9�n�9Yq�9!s�9�t�9�t�9�o�9�p�9u�9ss�9x   x   �v�9�u�9yr�9�q�9�o�9�s�9pr�9+p�9�o�9�q�9=r�9up�9Ks�9$p�9Aq�9.s�9�t�9�v�9�q�9.t�9�w�9�s�9=y�92t�9�s�9�x�9s�9�v�9+u�9r�9x   x   -u�9�s�9*p�9gp�9s�9Vt�9�o�9t�9Eq�9�q�9�o�9�u�92r�9Aq�9+p�9,s�9�v�9w�9�r�9�s�9c{�9x�9Iu�9�v�9�t�9&z�9�z�9t�9/r�9�v�9x   x   _y�9�r�9t�9�t�9�u�9�p�9p�9*t�9�t�93q�96p�9�u�9�t�9+s�9/s�9$y�9Yu�9nu�9�u�9�t�9Qy�9�u�93{�9�|�91t�9x�9�u�9�t�9v�9�v�9x   x   �v�9�s�9as�9~o�9zo�9u�9�t�9�p�9?t�9�t�9�n�9�o�9�s�9�t�9�v�9Uu�9jr�9�x�9x�9Lv�9�t�9x�9�z�9zx�9Fv�9Xv�9�w�9�y�9p�9u�9x   x   [w�9�u�9Pr�9rp�9Yp�9q�9sn�9pn�9�p�9|q�9q�9�q�9iu�9�v�9!w�9nu�9�x�9y�9�x�9�z�9Ay�9%~�9b|�9�x�9�y�9�x�9�x�9�y�9�w�9Nv�9x   x   ]q�9�m�9�o�9�t�9�p�92l�9�m�9$m�9`p�9Xs�9�o�9wn�9r�9�q�9�r�9�u�9x�9�x�9,z�9�|�9nz�9h}�9�|�9=|�9*{�9�y�9!w�9Gt�9�q�9pr�9x   x   �p�9-n�9�k�9o�9�l�9�s�9�r�9�l�9�p�9�l�9�m�9p�9St�9+t�9�s�9�t�9Nv�9�z�9�|�9w|�9�y�9�x�9�{�9C}�9�x�9sv�9�v�9Vt�9Cu�9�s�9x   x   *t�9�n�9�l�9�o�9�o�9[s�9�q�9n�9<k�9�n�9nu�9�p�9�u�9�w�9c{�9Oy�9�t�9>y�9nz�9�y�95{�9�y�9�z�9z�9v�9�w�9Yz�9�v�9�t�9�q�9x   x   Wr�9�o�9sk�9�n�9ij�9�h�9En�9�m�9gp�95q�9"n�9gp�9�n�9�s�9x�9�u�9x�9%~�9h}�9�x�9�y�9�}�9�|�9�v�9�u�9�y�9t�9p�9�p�9Nm�9x   x   �o�9�l�92m�9o�9�j�9"p�9�l�9j�9q�9�m�9t�9?v�9Wq�9:y�9Iu�9/{�9�z�9f|�9�|�9�{�9�z�9�|�9A}�9\{�9u�9	x�9�p�9#u�9�s�9�n�9x   x   Ui�9�i�9�o�9Bl�9�l�9o�9k�9 j�9Zm�9�p�9�r�9wo�9!s�93t�9�v�9�|�9yx�9�x�9;|�9>}�9$z�9�v�9]{�9!w�9�s�9�t�9�o�9�s�9�p�9�l�9x   x   �o�9�l�95m�9Kn�9�l�9ul�9Fo�9�k�9Ol�9�n�9�q�9wu�9�t�9�s�9�t�92t�9Bv�9z�9+{�9�x�9|v�9�u�9u�9�s�9�t�9"t�9Cq�9#m�9 l�9'n�9x   x   �k�9�g�9�h�9Wi�9Yi�9�i�9�k�9:s�99o�9�o�9�u�9�s�9�t�9�x�9$z�9x�9\v�9�x�9�y�9xv�9�w�9�y�9	x�9�t�9&t�9�v�9^p�9�q�9 q�9i�9x   x   �i�9ah�9<i�9�f�9Cj�9/h�9�i�9Jn�9�n�9]q�9r�9�o�9�o�9s�9�z�9�u�9�w�9�x�9w�9�v�9Xz�9t�9�p�9�o�9Gq�9bp�9	m�9�m�9�l�9bh�9x   x   j�9�h�9}j�9"j�9gj�9�n�97f�9�l�9so�9�l�9�s�9�u�9�p�9�v�9
t�9�t�9�y�9�y�9Dt�9Tt�9�v�9 p�9%u�9�s�9$m�9�q�9�m�9e�9m�9j�9x   x   !k�9�f�9"j�9�g�9�h�9�m�9Vk�9�r�9n�9Pp�9�s�9�o�9u�9,u�9-r�9v�9�o�9�w�9�q�9Ju�9�t�9�p�9�s�9�p�9�k�9"q�9m�9m�9aj�9_h�9x   x   �d�9d�9 f�9Tj�9,i�9�h�9.j�9�k�9�k�9�o�9�m�92r�9ws�9r�9�v�9�v�9u�9Jv�9kr�9�s�9�q�9Lm�9�n�9�l�9&n�9i�9kh�9j�9_h�9Td�9x   x   ;��9Ѧ�9ۤ�9��90��9&��9��9���9Ү�9G��9V��9S��9H��9ݳ�9��9���9g��9)��9��9��9ԯ�9���9��9ԭ�9K��9 ��9��9S��9q��9	��9x   x   Φ�99��9���91��9]��9b��9Z��9l��9p��9���9��9w��9z��9��9^��9���9=��9ѳ�9���9��9o��9���9��9e��9���9���9���9P��9���9z��9x   x   ؤ�9���9ɧ�9)��9��9@��9e��9A��9���9���9��9*��9��9n��9O��9-��9��9���9}��9��9Ӱ�9���92��9z��9A��9c��9��9���9@��9���9x   x   ��9/��9(��9���9��9���9ب�9��9���9ٯ�9���9X��9��9@��9���9���9���9���9 ��9���9ΰ�9 ��9���9���9H��99��9��9��9���9���9x   x   2��9Z��9��9��9���94��9ͫ�9���9���9L��9���9̮�9���9Ű�9��9��9���9��9���9���9��9���9��9���9���9��9!��9W��9u��9ʡ�9x   x   )��9a��9=��9���97��9_��9Ǩ�9ױ�9ݭ�9��9˰�9���9s��9z��9���9ۯ�9��9ϭ�9`��9Y��9=��9٬�9��9��9��9���9���9��9���9���9x   x   ��9W��9b��9٨�9ʫ�9Ǩ�9װ�9���9ԭ�9q��9~��9&��9���9D��9���9%��9���9@��9±�9���9��9q��9n��9���99��9<��9f��9
��9٧�9��9x   x   ���9l��9@��9��9���9ױ�9���9���9���9ų�9���9;��9M��99��9���9f��9���9���9���9���9!��9��9��9z��9֬�94��9֭�9G��9���9���9x   x   Ӯ�9p��9���9���9���9ܭ�9ԭ�9���9���9���9���9���9���9��9@��9-��9}��9��9���9���9���9���9���9ȯ�9���9���9r��9N��9̬�9L��9x   x   E��9���9���9ٯ�9H��9��9p��9���9���9]��9X��9R��9B��9��9C��9H��9���9 ��9r��9J��9��9���9���9l��9���9���9:��9V��9B��9ѭ�9x   x   Q��9��9��9���9���9Ȱ�9~��9���9��9V��9���9F��9��9m��9 ��9��9���9��9Z��9J��9q��9���9���9���9��9��9��9���9��9ʴ�9x   x   P��9y��9(��9_��9ͮ�9���9+��9:��9���9Q��9E��9��9���9���9Ѳ�9گ�9���9���9ִ�91��9k��9���9���9@��9Я�9r��9��9ί�9M��9ή�9x   x   F��9~��9��9��9���9q��9���9M��9���9F��9��9���9ǲ�9���97��9���9U��9p��9���9;��9���9*��98��9>��9���9!��9��9���93��9���9x   x   ׳�9��9m��9;��9���9w��9F��95��9��9���9h��9���9���9��9*��9��9,��9 ��9��9c��9���9���9ڷ�9w��9?��9���9��9��9���9y��9x   x   ��9`��9Q��9���9��9���9���9���9A��9E��9%��9Ҳ�96��9.��9���9��9(��9Q��9"��9
��9���9���9³�9h��9���9���9װ�9$��9��9���9x   x   ���9���9/��9���9 ��9ۯ�9)��9e��92��9J��9��9ޯ�9���9��9��9ܱ�9��9+��9N��9ƶ�9��9���9w��9%��9���9I��9ɷ�9��9q��9:��9x   x   j��9?��9��9���9���9��9���9���9}��9���9���9���9T��9,��9(��9��9$��9���9���9R��9���9���9r��9��9A��9c��9��9��9��9��9x   x   (��9ʳ�9���9���9��9̭�9C��9��9��9%��9��9���9g��9"��9U��9,��9���9���9\��9 ��9>��9���9��91��9ݸ�9p��9��9g��9��9���9x   x   ��9���9��9��9���9_��9ʱ�9���9���9o��9]��9մ�9���9��9!��9O��9���9U��9���9O��9���9%��9M��9Ӽ�9ȶ�9���9���9\��9 ��9ӳ�9x   x   ��9��9��9���9���9W��9���9���9���9G��9M��94��9?��9c��9��9Ƕ�9R��9���9P��9ϸ�9ü�9P��9��9޽�9��9޺�9,��9���9��9 ��9x   x   ӯ�9o��9ϰ�9Ͱ�9��9?��9��9��9���9��9r��9h��9���9���9���9��9���9A��9���9ü�9w��9ż�9��9��9Z��9���9���9��9o��9��9x   x   ���9���9��9#��9���9ج�9u��9��9���9���9���9���9+��9���9���9���9���9���9"��9Q��9Ƽ�9���9m��9ٹ�9ֻ�9o��9���9���9q��9
��9x   x   ��9��9-��9���9��9��9m��9��9���9���9���9���9>��9ַ�9���9z��9o��9��9L��9��9��9g��9��9ٷ�9��9Զ�9���9ӯ�9���9���9x   x   ڭ�9g��9t��9Ĥ�9���9��9���9��9Ư�9q��9���9D��9H��9u��9g��9%��9��94��9׼�9��9��9չ�9Է�9���9���9���9���9O��9���9���9x   x   J��9���9@��9G��9���9��9:��9ج�9���9���9��9ʯ�9���9=��9���9���9?��9ݸ�9Ͷ�9��9V��9ڻ�9��9���9��9e��9ݳ�9���9W��92��9x   x   ���9���9d��9<��9��9���9=��9:��9���9���9��9m��9'��9���9���9N��9_��9h��9���9޺�9���9o��9Ѷ�9���9f��9��9!��9Z��9M��9O��9x   x    ��9���9��9��9%��9���9h��9֭�9n��9:��9 ��9��9��9��9ٰ�9ͷ�9��9��9���90��9���9���9���9���9س�9 ��9h��9c��9���9���9x   x   Y��9Q��9���9 ��9]��9��9
��9L��9M��9W��9���9̯�9���9��9#��9��9��9d��9Z��9���9��9���9ү�9P��9���9\��9h��9֥�9J��9���9x   x   m��9���9@��9���9t��9���9է�9���9̬�9H��9��9Q��96��9���9��9|��9��9��9��9��9q��9v��9���9���9V��9G��9���9E��9��9��9x   x   
��9~��9���9���9ʡ�9���9��9���9L��9ͭ�9ʴ�9Ǯ�9���9z��9���9<��9��9���9ѳ�9���9ݭ�9��9���9���94��9M��9���9��9��9ª�9x   x   5��9���9R��9E��9���9��9P��9Q��9���9���9���9���9���92��9s��9���9H��9���9*��9���9/��9���9f��9M��9w��9���9��94��9���9���9x   x   ���9���9���9d��9���9���9=��9��9���9���9���9��9���9���9���92��9*��9��9���9���9���9s��9���9���9j��9���9���9���9!��9��9x   x   V��9���9>��9���9��92��9k��9��9���9���9���9���9���9;��9)��9��9k��9���9
��9���9���99��9C��9���9���9���9���9z��9l��9���9x   x   D��9b��9���9 ��9���9_��9���9���9���9>��9���9���9���9k��9'��9���9���9���9���9���9���9H��9���9��9���9��9��9:��9���9i��9x   x   ���9���9��9���9D��9X��9���9^��9l��9��9U��95��9`��9p��9���9j��9��9��9��9���9��9���9O��9���9G��9���9s��9���9w��9���9x   x   ��9���92��9_��9X��9���9E��9��9���9H��9���9���9��9K��9W��9���9?��9~��9���9s��9���9���9��9���94��9l��9G��90��9���9o��9x   x   N��9?��9i��9���9���9F��9]��9~��9��9���9���9���9���9j��9���9���9��9���9��9^��9��9���9���9��9���9���9���9���9\��9��9x   x   U��9��9��9���9_��9	��9���9���9q��9h��9��9���9���9���9F��9���9��9F��9���9��9���9��9���9���9���9���9���9���9���97��9x   x   ���9���9���9���9k��9���9��9u��9���9@��9���9q��9/��9{��9X��9���9���99��9���9���9���9Z��9E��9���9���9`��9��9���9<��9/��9x   x   ���9���9���9=��9��9H��9���9l��9?��9$��9v��9F��9���9���9l��9���9w��9l��9��9���9���9��9���9���9<��9"��9M��9��9���9���9x   x   ���9���9���9���9U��9���9���9��9���9q��9���9w��9���9,��9$��9���9���9���9t��9���9~��9���9O��9W��9���9%��9F��9���94��9%��9x   x   ���9��9���9���94��9���9|��9���9o��9D��9x��9���9l��9���9���9���9e��9���94��9���9���9A��9���9���9���9H��9 ��9"��9���9��9x   x   ���9���9���9���9d��9��9���9���9*��9���9���9k��9���9���9���9���9���9��9���9v��9���9@��9:��9W��9T��9W��9���9���9A��9���9x   x   /��9���98��9o��9w��9M��9i��9���9~��9���9-��9���9���9��9���9W��9���9<��98��9Y��9j��9c��92��9���9	��9,��9���9���9���9n��9x   x   s��9���9(��9,��9���9X��9���9H��9[��9i��9#��9���9���9���9���9���9��9���9��9f��9<��9���9���99��9���9���9���9���9;��9���9x   x   ���9.��9��9���9c��9���9���9���9���9���9���9���9���9V��9���9g��9���9��9���9���9���9��9&��9 ��9+��9���9���9���9]��9u��9x   x   E��9)��9n��9���9}��9B��9��9��9���9y��9���9e��9���9���9��9���9>��9���9��9:��9���9���9� �9���9J��9m��9���9n��9���9���9x   x   ���9��9���9���9��9{��9���9C��99��9m��9���9���9��9=��9���9��9���9���9���9V��9�9��9!�9��9���9���9%��9N��9-��9Q��9x   x   +��9���9
��9���9��9���9���9���9���9��9v��94��9���94��9��9���9��9���9��9���9���9'��9���9���9���9k��9���9e��9i��9���9x   x   ���9���9���9���9���9p��9^��9 ��9���9���9���9���9t��9_��9k��9���9@��9T��9���9( �9. �9� �9� �9
��9���9���9A��9���9m��9���9x   x   2��9���9���9���9��9���9 ��9���9���9���9���9���9���9f��9=��9���9���9�9���91 �9���92 �9(��92�9p��9��9���9���9���9j��9x   x   ���9x��9<��9H��9���9���9���9"��9^��9��9���9G��9B��9b��9���9��9���9��9&��9� �92 �9>��9A�9���9���9���9���9��9���9���9x   x   d��9���9G��9���9L��9��9��9���9G��9���9O��9���96��97��9���9)��9� �9#�9���9� �9'��9B�9@ �9q��9���9���9���9���9���9���9x   x   O��9���9���9��9���9���9��9���9���9���9U��9���9R��9���96��9��9���9��9���9��90�9���9m��9t��9[��9���9y��9@��9|��9��9x   x   x��9n��9���9���9I��94��9���9���9���99��9���9���9U��9��9���9+��9O��9���9���9���9r��9���9���9[��9���97��9T��9��9���9���9x   x   ���9���9���9��9���9n��9���9���9h��9!��9+��9L��9Q��93��9���9���9q��9���9n��9���9��9���9���9���99��9���9���9���9"��9���9x   x   ���9���9���9��9p��9G��9���9���9��9H��9M��9$��9���9���9���9���9���9)��9���9B��9���9���9���9��9V��9���9F��9��9j��9���9x   x   2��9���9~��98��9|��92��9���9���9���9��9���9&��9���9���9���9���9p��9Q��9f��9���9���9��9���9E��9��9���9��9W��9���9��9x   x   ���9��9k��9���9u��9���9\��9���9?��9���90��9���9?��9���9:��9\��9���9,��9g��9h��9���9���9���9��9���9#��9n��9���9x��9I��9x   x   ���9��9���9m��9���9s��9��9:��9/��9���9$��9��9���9m��9���9v��9���9S��9���9���9l��9���9���9��9���9���9���9��9J��9���9x   x   ."�9e$�9}%�90$�9�$�9c'�96+�9�,�9�4�94�9�3�98�9�8�9�8�9U9�9�:�9-9�9z7�9]9�9�7�94�94�95�9z-�9+�9'�9%�9�$�9�#�9E$�9x   x   b$�9�!�9�"�9#$�9�(�9`*�9�)�9�-�91�972�9N3�9�:�9�9�9n5�9n7�9m7�9S6�9�9�97;�93�9�1�9�1�9p,�92*�9�*�9q(�9�#�9�"�9�"�9z$�9x   x   {%�9�"�9u&�9�&�9'�9	)�9)+�9!.�9�/�9A1�9S5�9�6�9�4�9�8�9w:�98�9�4�9�5�9�5�9	2�9K/�9�.�9�+�9R(�9?'�9'�9Y&�9�"�9$�9r$�9x   x   0$�9&$�9�&�9�$�91*�9�*�9D/�9�0�9~4�9y8�9j4�9�0�997�98�99�9K7�9�1�9�4�9D7�9�4�9�0�9/�9+�9�*�9�#�9�&�98$�9�$�9�"�9� �9x   x   �$�9�(�9'�9-*�9:'�94(�9�.�9�.�9�2�9s2�9�1�9�7�9�6�9�1�9q6�97�91�9u3�9�2�9/�9�.�9�'�9"'�9�*�9�'�95(�9�$�9�%�9�!�9y&�9x   x   d'�9]*�9)�9�*�91(�9�.�9d1�990�9\3�9�1�9�5�9.5�9~3�9�2�9�6�9�6�9�0�9�3�90�9�0�9�.�9�(�9.*�9�(�9*�9�'�9�$�9�"�9l#�9$�9x   x   7+�9�)�9++�9E/�9�.�9e1�9�1�9�3�9G5�9	2�9�4�9 5�9�6�9�4�9�2�9+3�9.5�9�3�9�2�9H1�9�-�9�/�9�+�9�)�9�+�9N)�9\)�9)�9�(�9�*�9x   x   �,�9�-�9".�9�0�9�.�990�9�3�9�2�9B3�94�9�6�9@5�9�5�9�7�9�3�9�2�9/3�9E3�9�/�9|/�9�0�9�-�98-�9�,�9	+�9*.�9s)�9*�9%.�9r*�9x   x   �4�91�9�/�9}4�9�2�9^3�9E5�9D3�99�944�9'5�9>5�9D3�9)5�9�8�9�2�9m5�9�3�9h2�9t4�9�/�981�9[5�9-�9�+�9./�9�+�94/�9#+�9�-�9x   x   4�932�9A1�9x8�9t2�9�1�92�94�914�9G1�9�6�9m8�9�0�9^3�9=5�9�1�9�1�9�2�9W8�9�0�9c2�9s3�9i3�9 2�9X+�9�1�9�0�9�+�92�9�2�9x   x   �3�9L3�9V5�9j4�9�1�9�5�9�4�9�6�9)5�9�6�9'5�9�6�9 6�9P6�94�96�991�9z4�9�5�953�9%4�9�+�9�5�98�9�-�9�6�9.�9�7�9�5�9,�9x   x   8�9�:�9�6�9�0�9�7�9.5�9 5�9F5�9B5�9t8�9�6�9~4�9�5�9z5�9�5�98�91�9\6�9�:�9�7�9�6�9)4�9M:�9�5�9�5�9!6�9�5�9�:�9J4�9/6�9x   x   �8�9�9�9�4�9<7�9�6�93�9 7�9�5�9C3�9�0�9�5�9�5�9�6�93�906�9M7�9�4�9:�9�9�9C8�9/<�98�9X6�9B:�9�;�9�9�9p6�9T7�9�<�9�8�9x   x   �8�9l5�9�8�98�9�1�9�2�9�4�98�9%5�9]3�9S6�9x5�93�932�9l8�9�8�9�5�9�7�9�9�9�<�9>>�9G;�9<�9w=�9�=�9�<�9r;�9�>�9�;�9�9�9x   x   R9�9m7�9v:�9�8�9n6�9�6�9�2�9�3�9�8�9?5�94�9�5�9/6�9g8�9g:�9�7�9�9�9�:�9�:�9n=�9�=�9�=�9�>�9�>�9">�9�<�9=>�9�=�9";�9�:�9x   x   �:�9r7�98�9P7�97�9�6�9(3�9�2�9�2�9�1�96�98�9Q7�9�8�9�7�9 :�9�9�9:�9'=�9#?�9�=�9�<�97@�9@�9�=�98>�9r>�9C=�9 :�9�9�9x   x   .9�9O6�9�4�9�1�91�9�0�9.5�923�9n5�9�1�9:1�91�9�4�9�5�9�9�9�9�9�:�9iC�9�?�9�B�9�A�99@�9�@�9�?�9�@�9�B�9b@�9�B�9l;�9�9�9x   x   y7�9�9�9�5�9�4�9t3�9�3�9�3�9G3�9�3�9�2�9z4�9U6�9:�9�7�9�:�9	:�9iC�9�?�9>?�9[C�9�A�9x@�9�@�9�A�9�C�9?�9�?�9�C�9Z9�9E;�9x   x   a9�93;�9�5�9D7�9�2�90�9�2�9�/�9e2�9X8�9�5�9�:�9�9�9�9�9�:�9'=�9�?�9>?�9 D�9�B�9�C�9�A�9*C�9C�9�C�9�>�9�?�9Y=�9;�9:�9x   x   �7�93�92�9�4�9/�9�0�9I1�9~/�9v4�91�993�9�7�9C8�9�<�9m=�9!?�9�B�9ZC�9�B�9�F�9 F�9eF�9�F�9mB�9eD�9�B�9�>�9�=�9�;�9}8�9x   x   4�9�1�9L/�9�0�9 /�9�.�9�-�9�0�9�/�9`2�9'4�9�6�9/<�9>>�9�=�9�=�9�A�9�A�9�C�9F�9lD�9�E�9D�9EA�9l@�9">�9>�9�>�9�<�9�6�9x   x   4�9�1�9�.�9
/�9�'�9�(�9�/�9�-�941�9k3�9�+�9(4�9 8�9L;�9�=�9�<�9:@�9v@�9�A�9_F�9�E�9�A�9�@�9�@�92=�9�=�9�:�9X7�9�3�9,�9x   x   
5�9m,�9�+�9+�9#'�9-*�9�+�9<-�9]5�9m3�9�5�9L:�9Y6�9<�9�>�99@�9�@�9�@�9/C�9�F�9D�9�@�9�?�98@�9�=�9�<�97�9�:�9}6�9l2�9x   x   v-�9.*�9V(�9�*�9�*�9�(�9�)�9�,�9-�92�9 8�9�5�9@:�9w=�9�>�9@�9�?�9�A�9C�9rB�9CA�9�@�94@�9c?�9�=�99�9�5�9M7�9&2�9�-�9x   x   +�9�*�9='�9�#�9�'�9*�9�+�9
+�9�+�9Y+�9�-�9�5�9�;�9�=�9">�9�=�9�@�9�C�9�C�9gD�9j@�9/=�9�=�9�=�96<�9I6�9X.�9�+�9�+�9�)�9x   x    '�9m(�9'�9�&�95(�9�'�9O)�9'.�91/�9�1�9�6�9!6�9�9�9�<�9�<�98>�9�B�9?�9�>�9�B�9">�9�=�9�<�99�9G6�9�5�9z1�9R.�9/�9�*�9x   x   %�9�#�9W&�95$�9�$�9�$�9a)�9w)�9�+�9�0�9.�9�5�9r6�9q;�9@>�9s>�9_@�9�?�9�?�9�>�9>�9�:�97�9�5�9W.�9�1�9P,�9�)�9�'�9g$�9x   x   �$�9�"�9�"�9�$�9�%�9�"�9)�9*�96/�9�+�9�7�9�:�9U7�9�>�9�=�9F=�9�B�9�C�9[=�9�=�9�>�9V7�9�:�9G7�9�+�9Q.�9�)�9�)�9�#�9&�9x   x   �#�9�"�9$�9�"�9�!�9j#�9�(�9#.�9"+�9!2�9�5�9I4�9�<�9�;�9";�9�9�9m;�9W9�9;�9�;�9�<�9�3�9~6�9&2�9�+�9/�9�'�9�#�9%!�9"�9x   x   D$�9{$�9q$�9� �9x&�9$�9�*�9p*�9�-�9�2�9,�936�9�8�9�9�9�:�9�9�9�9�9E;�9:�9�8�9�6�9,�9n2�9�-�9�)�9�*�9d$�9�%�9�!�9%�9x   x   0c�9�^�9 c�96a�9i�9�h�9�h�9�p�9m�9�r�9n}�9jy�9�|�9�~�9v�9��9"~�9C~�9�|�9�x�9�}�9{q�9�m�9�q�9�i�9�h�9�g�9�a�9�`�9�^�9x   x   �^�9�[�9�d�9d�9Oh�9Zh�9�k�9�r�9"p�9t�9�x�91v�9j{�9�|�9�|�9�}�9�}�9�z�9�v�9Mx�9�t�9sq�93p�9�k�9�g�9�h�9hd�9qf�9	]�9�]�9x   x   �b�9�d�9yf�9�e�9Qg�9lm�9�k�9�q�9t�9�t�9�w�9sx�9 |�9k}�9�|�9Z|�9�{�9Yx�9 x�9St�9Ar�9�r�9m�9�l�9bg�9�f�9Jd�9d�9Yc�9mg�9x   x   5a�9d�9�e�9�h�9~j�9�p�9�k�9@r�9Lt�9	r�9�{�9n|�9�x�9�{�9�|�9Wy�9�}�9.z�9Er�9v�9r�9k�9no�9�k�9�f�9g�9
f�9�`�9\c�9~b�9x   x   i�9Ph�9Tg�9j�9vm�9Cu�9p�9u�9|r�9Mu�9�{�9!z�99y�9�{�9y�9�x�9�{�9�v�9p�9Fu�9�p�9Nu�9bm�9k�9�g�9�f�9�h�9�e�9�f�9�f�9x   x   �h�9Yh�9km�9�p�9Cu�9�p�9Vn�9[s�9�u�9�x�9x�9�x�90|�9l{�9`z�9qx�9�w�9�v�9�t�9Em�9�p�9�v�9�n�9�m�9�h�9�h�9ll�9�m�9Ym�9k�9x   x   �h�9�k�9�k�9�k�9p�9Sn�9�v�9.x�9�u�9�y�9�y�9�x�9az�9^x�9�x�9�z�9�t�9�w�9�v�9_o�9n�9l�9�l�9vj�9ej�9>h�9�g�9#j�9�h�9�i�9x   x   �p�9�r�9�q�9;r�9u�9[s�9-x�9Hr�9u�9]y�9�w�9x�9My�9]x�9�x�9�u�9�r�9�w�9Es�9�u�9*s�92q�9�r�9#p�9�p�9.n�9o�9�n�9�l�9�p�9x   x   m�9p�9 t�9Mt�9|r�9�u�9�u�9u�9Cy�9�x�9]x�9�w�9'w�9�y�97x�9Vt�9
v�9�v�9�p�9At�9�s�9�o�9wn�9\p�9�p�9]r�9�p�9s�9�p�9�p�9x   x   �r�9�s�9�t�9r�9Iu�9�x�9�y�9[y�9�x�9{z�9 y�9?z�9�y�9�x�9{�9�y�9�w�9v�9os�9�s�9�u�9�q�9�s�9�t�9ou�95r�9:q�9{v�9t�9t�9x   x   l}�9�x�9�w�9�{�9�{�9x�9�y�9�w�9]x�9y�9w�99y�9�x�9!w�9Kx�9�y�9�{�9Zz�9:w�9�x�9�|�9�y�9_w�9Pw�9�|�9}�9�{�9{v�9w�9�y�9x   x   ky�91v�9vx�9n|�9#z�9�x�9�x�9wx�9�w�99z�93y�9Qw�9�x�9z�9�x�9�x�9j}�9�x�9�v�9�x�9�y�9|�9�w�9�w�9�v�9-x�9�x�9y�9�{�9�x�9x   x   �|�9f{�9�{�9�x�99y�91|�9_z�9Hy�9)w�9�y�9�x�9�x�9;y�9�{�9�y�9y�9w{�9�z�9�|�9�x�9�{�9 }�9���9���9�z�9�~�9��9�{�9�}�9�x�9x   x   �~�9�|�9i}�9�{�9�{�9o{�9]x�9Zx�9�y�9�x�9w�9z�9�{�9�{�9
|�9�|�9�}�9�~�9\}�9���9��9T��9q��9���9���9M��9��9��9@�9}�9x   x   y�9�|�9�|�9�|�9y�9bz�9�x�9�x�99x�9{�9Jx�9�x�9�y�9|�9}�9 }�9�~�9��9Ѐ�9H�9��9��9���9���9d��9�~�9g��9�9V��9*��9x   x   ��9�}�9Z|�9Sy�9�x�9sx�9�z�9�u�9[t�9�y�9�y�9�x�9y�9�|�9!}�9���9^��9��9��9���9���9ʉ�9؉�9���9ڋ�9!��9��9U��9���9���9x   x   #~�9�}�9�{�9�}�9�{�9�w�9�t�9�r�9v�9�w�9�{�9i}�9{{�9�}�9�~�9Y��9 ~�99��9L��9A��9���9��9$��9���9���9���9Ȇ�9��9{��9���9x   x   F~�9�z�9]x�9.z�9�v�9�v�9�w�9�w�9�v�9v�9]z�9�x�9�z�9�~�9��9��95��9c��9��9��9���9���9��9g��9]��9$��9���9��9��9���9x   x   �|�9�v�9�w�9Ar�9p�9�t�9�v�9Ds�9�p�9ns�98w�9 w�9�|�9`}�9π�9$��9J��9!��9͌�9+��9��9��9 ��9t��9���9���9Ά�9��9	��9S}�9x   x   �x�9Ox�9Vt�9v�9Cu�9Hm�9ao�9�u�9At�9�s�9�x�9�x�9�x�9���9F�9���9?��9
��9-��9o��9���9���9B��9���9/��9��9���9^�9�~�9y�9x   x   �}�9�t�9>r�9r�9�p�9�p�9n�9.s�9�s�9�u�9�|�9�y�9�{�9��9��9���9���9���9��9���9���9���9�9��9���9��9��9~��9'}�9�y�9x   x   �q�9uq�9�r�9k�9Ou�9�v�9	l�93q�9�o�9�q�9�y�9|�9 }�9P��9��9Ή�9��9���9��9���9���9Ŏ�9���9��9���9��9 ��9V|�9�z�9ty�9x   x   �m�97p�9}m�9po�9dm�9�n�9�l�9�r�9vn�9�s�9aw�9�w�9���9p��9���9؉�9#��9��9��9=��9���9���9��9���9���9��9ـ�9jx�97y�9�s�9x   x   �q�9�k�9�l�9�k�9 k�9�m�9xj�9&p�9Xp�9�t�9Ow�9x�9���9���9���9���9���9h��9t��9���9��9��9���9Ҁ�9M��9�~�9:x�9v�9Gs�9�p�9x   x   �i�9�g�9dg�9�f�9�g�9�h�9fj�9�p�9�p�9ru�9|�9�v�9�z�9���9c��9ߋ�9���9\��9���9-��9���9���9���9L��9�z�9Cx�9�|�9dv�9�q�9�n�9x   x   �h�9�h�9�f�9g�9�f�9�h�9>h�92n�9Xr�9<r�9}�9-x�9�~�9J��9�~�9(��9݆�9-��9���9��9��9��9��9�~�9Fx�9�z�9�r�9�p�9�n�9�i�9x   x   �g�9kd�9Nd�9f�9�h�9jl�9�g�9o�9�p�9Bq�9�{�9�x�9��9��9g��9��9Ɔ�9���9ӆ�9���9��9"��9ـ�99x�9�|�9�r�9�p�9qo�9�f�9Sl�9x   x   �a�9qf�9d�9�`�9�e�9�m�9j�9�n�9s�9|v�9|v�9y�9�{�9��9�9[��9��9��9���9[�9~��9X|�9lx�9v�9dv�9�p�9oo�9�j�9�m�9�f�9x   x   �`�9]�9Yc�9Vc�9�f�9Zm�9�h�9�l�9�p�9t�9�w�9�{�9�}�9>�9W��9���9|��9��9��9�~�9$}�9�z�99y�9Is�9�q�9�n�9�f�9�m�9	f�9�b�9x   x   �^�9�]�9ng�9{b�9�f�9k�9�i�9�p�9�p�9t�9�y�9�x�9�x�9}�9/��9��9���9���9R}�9y�9�y�9ry�9�s�9�p�9�n�9�i�9Tl�9�f�9�b�9di�9x   x   l��9���9���9Ҧ�9��9���9���9���9)��9���9и�9���9���9���9��9���9 ��93��9���9ھ�9k��9���9ҳ�9���9E��9���9z��9i��9��9X��9x   x   ���9%��9z��9���9n��9���9ΰ�9��9���9!��9\��9Ͻ�9���9���9���9���9���9˿�9{��9=��9���9%��9S��9���9���9��9إ�90��9��9���9x   x   ���9}��9x��9c��9v��9K��9���9���9��9Z��96��9i��9>��9d��9ؽ�9n��9L��9a��9���9���9k��9T��9&��9"��9z��9��9@��95��9��9��9x   x   Ц�9���9^��9���9w��9��96��9ǲ�9���9m��9���9̾�9^��9о�9*��9��9п�9q��9+��9q��9���9���9ȭ�9Ь�9H��9���9��9J��99��9���9x   x   ��9r��9u��9y��9M��9̮�9<��90��9���9:��9.��9��9��9u��9��9���9��9r��9���9d��93��9\��9��9���9��9O��9���9΢�9
��91��9x   x   ���9���9G��9��9Ǯ�9��9_��9v��9���9���9T��9��9���9��9��95��9׻�9ü�9g��9|��9ر�9��9���9���9\��9���9ܧ�9K��9��9��9x   x   ���9а�9���99��9=��9Y��9?��9s��9��9^��9���9���9��9��9���9���9 ��9L��9߶�9>��9��9��9���9ܮ�9Ȯ�9���9���9��9O��9��9x   x   ���9��9���9Ʋ�95��9v��9t��9���9���9��9��9D��9���9���9��9���9;��9\��9���9=��9���9M��9��9��9-��9@��9��9	��9��9��9x   x   ��9���9��9���9���9���9��9���9���9���9(��9���9-��9���9��9���96��99��9���9ݴ�9���9��9%��9���9��9Ǳ�9��9���9N��9��9x   x   ���9&��9Y��9q��9?��9���9b��9��9���9���9��9Y��9��9��9ּ�9���9Y��9���9��9��9Ժ�9��9G��9*��9ڹ�9��9���9#��9���9p��9x   x   ָ�9^��9/��9���9/��9N��9���9��9*��9��9ܼ�9*��9l��9��9���9���9?��9���9��9���9p��9D��9���9��9H��9ε�9x��9���9��9���9x   x   ���9ҽ�9i��9Ǿ�9��9��9���9G��9���9Z��9'��9���9S��9M��9S��9G��9Q��9j��9��9˿�9���9���9s��9���9���9���9���9��9���9���9x   x   ���9���9>��9\��9��9���9��9���9.��9��9l��9S��9b��9N��9&��9s��9^��9_��9���9���9���9���9.��9���9���9	��9j��9f��9Z��9���9x   x   ��9���9f��9ξ�9u��9���9	��9���9���9��9��9O��9G��9��9���9���9~��9Z��9���9���9k��9���9p��9���9b��9���9���9��9n��9���9x   x   ��9���9Խ�9+��9��9��9���9��9��9Ѽ�9���9X��9(��9���9`��9���9���9J��9C��9���93��9S��9Z��9S��9��9/��9&��9���9-��9���9x   x   ���9���9m��9��9���91��9���9���9���9���9���9F��9s��9���9���9���9���9���9���9���9���9��9���9��9���9��9���9G��9%��9l��9x   x   ���9���9L��9ο�9��9ػ�9��9@��98��9^��9D��9P��9\��9���9���9���9���9��9���9u��9���9���9?��9���9���9���9���9���9@��9|��9x   x   2��9Ͽ�9c��9q��9u��9���9R��9a��97��9���9���9n��9^��9^��9M��9���9��9���9���9���9���9"��9M��9x��9���9\��9���9<��9,��9��9x   x   ���9|��9���9,��9���9e��9ݶ�9���9ü�9��9}��9��9���9���9A��9���9���9���9���9���9���9���9���9���9	��9l��9���9���9:��9O��9x   x   ھ�9=��9���9p��9c��9}��9@��9:��9��9��9���9п�9���9���9~��9���9w��9���9���95��9���9���9���9���9���9���9��9T��9���9���9x   x   j��9���9m��9���91��9۱�9��9���9���9Ӻ�9k��9���9���9p��93��9���9���9���9���9���9=��9���9��9H��9��9���9���9n��9���91��9x   x   ���9%��9V��9���9\��9��9��9O��9��9��9@��9���9���9���9Y��9
��9���9'��9���9���9���9���9���9���9d��9|��9���9C��9��9���9x   x   ɳ�9V��9'��9ʭ�9��9���9���9��9#��9H��9���9{��9,��9t��9_��9���9?��9K��9���9���9��9���9���9���9h��9���9>��9���9ع�9T��9x   x   ���9���9 ��9Ь�9���9���9ۮ�9��9���9-��9��9���9���9���9V��9��9���9|��9���9���9K��9���9���9���9+��9A��9���9P��9���9��9x   x   C��9���9z��9H��9��9b��9Ʈ�9,��9��9ݹ�9J��9���9���9e��9��9���9���9���9��9���9��9^��9e��9+��9���9[��9��9&��9���9c��9x   x   ���9��9��9���9O��9��9���9A��9ɱ�9��9ѵ�9���9	��9���93��9��9���9_��9h��9���9���9x��9���9D��9[��9(��98��9���9>��9-��9x   x   x��9ץ�9>��9��9���9ާ�9���9%��9��9���9{��9���9f��9���9%��9���9���9���9���9��9���9���9=��9���9��92��9I��9T��9/��9/��9x   x   g��90��92��9L��9ˢ�9O��9��9��9���9$��9���9��9j��9��9���9I��9���9:��9���9Y��9p��9D��9���9V��9'��9���9W��9��9n��9Z��9x   x   ���9���9��9<��9
��9��9N��9��9O��9���9��9���9Y��9s��9+��9"��9E��9)��9;��9���9���9��9Թ�9���9���9;��9-��9o��9+��9��9x   x   Y��9���9���9���9-��9��9��9��9��9o��9���9���9���9���9���9k��9y��9���9P��9���90��9���9U��9��9b��9+��9,��9[��9��9��9x   x   ���9��9v��9���91��9S��9��9��9���9Z�9��9D�99�9A
�9��9��9��9D�9��9-�9�92��9H��9��9���9��9 ��9`��9}��9���9x   x   ��9���9���96��9N��9���97��9���9k��9���9W �9H
�9T
�9a�9�9��9��9��9[
�9I�9( �9���9���9��9��9���9���9���9"��9���9x   x   s��9���9U��9B��9���9B��9���9E��9���9� �9��9{�9��9�
�9��9�	�9��9��9��9*��9���9���97��9\��9*��9���9��9���9���9���9x   x   ���97��9B��9 ��9���9���9���96��9���9�9��9N�9��9,�9\�9b�9��9��9�9���9A��9���9#��9���9���9���9��9/��9_��9���9x   x   /��9M��9���9���9��9���9���9U��9���97 �9`�9
�9��9B�9��98	�9��9	�9���9���9$��9I��9J��9���9���9���9<��9!��9���9H��9x   x   R��9���9D��9���9���9Q��95��9���9Y �9��9��9M�9�9x�9��9��9s�9� �9Y��9���9���9���9���9b��9&��9 ��9���9���9@��9��9x   x    ��95��9���9���9���91��9� �9��9���9>�9��9��9��9T�9r�9)�9&��9��9y��9��9���9z��9Q��9P��9���9���9���9��9���9��9x   x   }��9���9A��95��9Z��9���9��9@ �9���9��9��9r�9J�9��9��9���9V �9��9���9���9���9g��9���9��9���9���9D��9	��9
��9a��9x   x   ���9m��9���9���9}��9Y �9���9���9��9��9��9K�9��9_�9]�9E��9���9��91��9q��9���9���98��98��90��9���98��9���9[��9���9x   x   Y�9���9� �9
�96 �9��9A�9��9��9� �9�9h�9���9��9.�9��9���9I �9��9���9���9D�9���9i��9k��9��9)�9u��9��9G��9x   x   ��9R �9��9��9`�9��9��9��9��9�9m
�9�9I�9��9��9��9��9)�9M�9� �9;�9w��9?�9��99��9^�9��9��9��9���9x   x   B�9J
�9{�9M�9
�9O�9��9q�9F�9l�9&�9�9T�99�9��9&�9��9��9 �9��9c�9.�9W
�9!�9��9��9r�9�	�9��9Y�9x   x   8�9N
�9��9��9��9�9��9E�9��9���9H�9N�9X�9��9D	�9��9��9��9��9��9��9��92�9��9��9�9��9��90�9w�9x   x   D
�9^�9�
�9(�9B�9w�9T�9��9_�9��9��98�9��9]�9��9Y
�9��9��9�
�9��9�9��9A�9Y�96�9��9��95�9��9�9x   x   ��9�9��9X�9��9��9u�9��9a�91�9��9��9C	�9��9P�9�
�9��9��9��9��9��9�9	�9U�9<�9��9f�9��9M�9�9x   x   ��9��9�	�9g�9?	�9��9(�9���9F��9��9��9)�9��9]
�9�
�9�9�9��9��9��9��9��9'�9��9��9�9��9��9$�9��9x   x   ��9��9��9��9��9v�9(��9T �9���9���9��9��9��9��9��9�9	�9$�9��9��9?"�9 �9#�9��9�!�9��9��9��9��9!�9x   x   E�9��9��9��9�9� �9��9��9��9D �9)�9��9��9��9��9��9&�9L�9 �9.!�9V�9X�9�9�9"�9��98�9b�9��9"�9x   x   ��9Y
�9��9�9���9a��9x��9���96��9��9Q�9 �9��9�
�9��9��9��9�9Y�9��9� �9��9��9��9-�9x�9��9f�9��93
�9x   x   2�9F�9+��9���9���9���9��9���9l��9���9� �9��9��9��9��9��9��9+!�9��9� �9�#�9�#�9�"�9F�9v"�9��9Y�97�9"�9��9x   x   �9' �9���9B��9#��9���9���9���9���9���9C�9j�9��9�9��9��9F"�9V�9� �9�#�9h�9�#�9?�9��9� �9��9 �9��9G�9��9x   x   3��9���9���9~��9K��9���9u��9k��9���9I�9u��90�9��9��9�9��9 �9T�9  �9�#�9�#�9X �9��9Q!�9L�93�9��9�9y�9���9x   x   N��9���98��9$��9K��9���9T��9���9:��9���9=�9Z
�93�9A�9�9+�9#�9�9��9~"�9@�9��9l �9f�9J�9��9��9�
�9��9S��9x   x   ��9��9]��9���9���9a��9S��9#��99��9l��9��9%�9��9Z�9U�9��9��9�9��9G�9��9M!�9g�9��9p�9�
�9�9�9U��9���9x   x   ���9��9'��9���9���9"��9���9���9-��9l��9>��9��9��97�9;�9��9�!�9"�9.�9y"�9� �9K�9O�9n�9��9�9���9���9���9L��9x   x   ��9���9���9���9���9��9���9���9���9��9]�9��9�9��9��9�9�9��9{�9��9��96�9��9�
�9{�9��9o�9���9w��9��9x   x   ���9���9	��9��9<��9���9���9A��9=��9(�9��9w�9��9��9i�9��9��94�9��9Y�9 �9��9��9�9���9p�9��9j��9���9)��9x   x   a��9���9���96��9"��9���9��9��9���9x��9��9�	�9��91�9��9��9��9b�9f�95�9��9�9�
�9�9���9���9k��9M��9���9[��9x   x   w��9 ��9���9b��9���9B��9���9
��9^��9��9��9��9/�9��9P�9"�9��9��9��9!�9K�9|�9��9V��9���9v��9���9���9z��9q��9x   x   ���9���9���9���9F��9��9��9b��9���9J��9���9]�9v�9�9�9��9"�9%�94
�9��9��9���9O��9���9M��9��9&��9U��9q��9��9x   x   ��9�"�9a%�99%�9(�9n0�9d4�9�;�9�=�9�D�9�N�9N�9yR�9MX�9�V�9�X�94U�9�X�9vS�9bM�9jN�9lC�9>�9>�9O3�9�/�9�(�9c%�9%�9�"�9x   x   �"�9"�9%*�9D&�9�+�9�/�9L7�9?=�9u=�93H�9&I�9�J�9LU�9�U�9T�9�T�9�V�90T�9'J�9DJ�9�H�9�=�9�;�9�6�91�9l,�9T%�9*�9�"�9�"�9x   x   c%�9#*�9�)�9�*�9�4�9r5�9i:�9�=�9`C�9yF�9H�9"L�9SS�9�S�9lN�9&S�9�R�9!M�9�G�9 E�9�C�9�>�9;�9r5�9/3�9�*�9�*�9�)�9
%�9�(�9x   x   >%�9D&�9�*�9W.�9�2�9�3�976�9A�9�E�9�F�9#Q�9�M�9	N�95M�9RM�96N�99N�9YP�9�G�9G�9�?�9�5�9h3�9�2�9|/�9p*�9�%�9u%�9�"�9O"�9x   x   (�9�+�9�4�9�2�9�3�9�9�9�<�93E�9<F�9	F�9"M�9L�9�N�9uP�9�N�9�K�9�L�9�F�9�D�9dE�9f>�9�9�9`3�92�9�3�9�+�9�(�9B*�9�%�9V*�9x   x   r0�9�/�9r5�9�3�9�9�9�B�9�A�9�E�9SI�9�J�9TJ�9J�9,R�9hQ�92J�9.K�9MJ�9rI�9�F�9�@�9�A�9]:�9�3�9�5�9�0�9]0�9r-�9Y,�9b,�9^.�9x   x   f4�9L7�9k:�986�9�<�9�A�9�C�9F�9�L�9�N�9�K�9nL�9/O�9M�9�J�9�N�9�L�9F�9�C�9aB�9=�9�5�9	;�9S6�9R3�9u0�9�+�9<0�9�*�9�/�9x   x   �;�9;=�9�=�9
A�92E�9�E�9F�9�E�9�L�9$K�9�L�9 L�9�K�9�L�9bK�9M�9�E�9�E�9�E�9 E�9MA�9?=�9d=�9&=�9�9�9E8�9�6�9�7�99�9e9�9x   x   �=�9t=�9cC�9�E�9;F�9WI�9�L�9�L�9�N�9J�9O�9�N�9�N�9�J�9�M�9PL�9qM�9�I�9�E�9�E�9D�9�=�9�<�9�<�9�?�9u?�9,7�9�>�9�?�9�=�9x   x   �D�9-H�9|F�9�F�9F�9�J�9�N�9%K�9J�9:O�91M�9 N�9N�9�I�9yL�9RN�9�I�9XF�9 H�9�E�9�G�9E�9B�95C�9�A�9�@�9�@�9)B�9vB�9�A�9x   x   �N�9'I�9H�9Q�9"M�9UJ�9�K�9�L�9O�91M�9�B�9OM�9P�9�K�9�J�9�K�9�M�9|O�9�G�9 J�99N�9�M�9mL�9�J�9�I�9�O�9J�9<K�9�L�9MM�9x   x   N�9�J�9#L�9�M�9L�9J�9nL�9%L�9�N�9�M�9NM�9N�9L�9�M�9�I�9_J�9O�9M�9^J�9�M�9Q�9cO�9�I�9�N�9P�9�O�9�M�9.I�9�O�93Q�9x   x   uR�9FU�9RS�9N�9�N�9*R�9-O�9�K�9�N�9�N�9P�9L�9�N�9�Q�9�O�9"N�9IR�9�T�9`R�9`Q�9�V�9xT�9tV�9�Y�9^R�9<Z�9�W�9T�9�V�9�P�9x   x   RX�9�U�9�S�9<M�9{P�9oQ�9M�9�L�9�J�9�I�9�K�9�M�9�Q�9�O�9�L�9�S�9�V�96Y�9�X�9�X�9n\�9V^�9 _�9V\�9�[�9^�9*^�9�\�9 Y�9RY�9x   x   W�9T�9iN�9TM�9�N�91J�9�J�9_K�9�M�9vL�9�J�9�I�9�O�9�L�9�N�9�S�9WU�9�Y�9�\�9]�9+_�9�_�9�^�9a�9�_�9�_�9l_�90\�9\�9�Y�9x   x   �X�9�T�9!S�93N�9�K�9,K�9�N�9M�9RL�9RN�9�K�9ZJ�9!N�9�S�9�S�9Z�9�Z�9i\�9�a�9�b�9�e�9f�9-f�9We�9�e�9�e�9c�9�b�9�\�9�Y�9x   x   4U�9�V�9�R�98N�9�L�9QJ�9�L�9�E�9pM�9�I�9�M�9O�9MR�9�V�9UU�9�Z�9�Y�9�`�9e�9�c�9d�9�g�9Hh�9�g�9Vd�9�c�9�d�9`�9�Z�9 \�9x   x   �X�91T�9)M�9VP�9�F�9wI�9F�9�E�9�I�9]F�9}O�9M�9�T�95Y�9�Y�9i\�9�`�9�g�9�k�9�e�9sh�9<l�9�l�9 h�9'f�9@l�9�h�9�`�9�Z�9Z�9x   x   xS�9%J�9�G�9�G�9�D�9�F�9�C�9�E�9�E�9$H�9�G�9bJ�9dR�9�X�9�\�9�a�9e�9�k�9�q�9�p�9*r�9�t�9�q�9�p�9Aq�9�j�9�d�9�c�9�\�9!X�9x   x   _M�9CJ�9 E�9G�9`E�9�@�9`B�9 E�9�E�9�E�9�I�9�M�9]Q�9�X�9]�9�b�9�c�9�e�9�p�9Am�9�o�90o�9n�9�p�9�f�9�d�9"a�9t\�9Y�9Q�9x   x   hN�9�H�9�C�9�?�9l>�9�A�9=�9XA�9D�9�G�97N�9Q�9�V�9m\�9,_�9�e�9d�9qh�9'r�9�o�9q�9�o�9Qq�9�g�9�b�91g�9%`�9
\�9W�9�P�9x   x   mC�9�=�9�>�9�5�9�9�9^:�9�5�9A=�9�=�9
E�9�M�9gO�9~T�9U^�9�_�9f�9�g�9=l�9�t�93o�9�o�9�t�91m�9Ei�9&e�9x^�9�^�9�S�9�O�99N�9x   x   >�9�;�9!;�9g3�9]3�9�3�9
;�9e=�9�<�9B�9oL�9�I�9zV�9!_�9�^�9.f�9Hh�9�l�9�q�9n�9Rq�97m�9�e�9�f�9$`�9�^�9�V�9�I�9�K�9"C�9x   x   >�9�6�9v5�9�2�92�9�5�9U6�9$=�9�<�97C�9�J�9�N�9�Y�9Y\�9a�9Ue�9�g�9h�9�p�9�p�9�g�9Ji�9�f�9g_�9E\�9�Y�9�N�9}K�9�B�9�;�9x   x   W3�9#1�9.3�9z/�9�3�9�0�9U3�9�9�9�?�9�A�9�I�9 P�9aR�9�[�9�_�9�e�9Yd�9(f�9@q�9�f�9�b�9)e�9"`�9C\�9�R�9�O�9�H�9�B�9�@�9�8�9x   x   �/�9o,�9�*�9m*�9�+�9^0�9t0�9K8�9x?�9�@�9�O�9�O�9BZ�9^�9�_�9�e�9�c�9Gl�9�j�9�d�9.g�9w^�9�^�9�Y�9�O�9EQ�9@�9G=�9P9�91�9x   x   �(�9R%�9�*�9�%�9�(�9p-�9�+�9�6�9.7�9�@�9J�9�M�9�W�9+^�9r_�9c�9�d�9�h�9e�9a�9*`�9�^�9�V�9�N�9�H�9@�9�9�9�6�9V*�9�-�9x   x   f%�9	*�9�)�9t%�9C*�9X,�9C0�9�7�9�>�9(B�99K�9,I�9T�9�\�9-\�9�b�9`�9�`�9�c�9u\�9\�9�S�9�I�9wK�9�B�9C=�9�6�9�0�9�,�9Q*�9x   x   %�9�"�9	%�9�"�9�%�9a,�9�*�99�9�?�9|B�9�L�9�O�9�V�9Y�9\�9�\�9�Z�9�Z�9�\�9�X�9	W�9�O�9�K�9�B�9�@�9P9�9W*�9�,�9K%�9�"�9x   x   �"�9�"�9�(�9P"�9_*�9].�9�/�9j9�9�=�9�A�9NM�97Q�9�P�9VY�9�Y�9�Y�9�[�9Z�9"X�9Q�9�P�96N�9&C�9�;�9�8�91�9�-�9T*�9�"�9�(�9x   x   �k�9�_�9kb�9�i�9Zl�9�s�9*{�9�{�9l��9��9��9ۗ�9���96��9��9���9���9��9j��9��9��9��9Q��9�|�9Tz�9�r�9�l�9mi�9d�9�_�9x   x   �_�9"b�9�e�9|i�9o�9�o�9�x�9��9��9;��9t��9���9���9��9D��93��9���9O��9|��9A��9��9���9Q�9x�9Jq�9)o�9ni�9�d�9a�9�_�9x   x   jb�9�e�9>c�9�m�9�r�9Zw�9�~�9x��9���9̐�9Ә�9G��9���9���9���9?��9���9R��9k��9G��9��9x��9��9w�9�q�9ym�9d�95f�9vc�96^�9x   x   �i�9xi�9�m�9�o�9Yt�9�}�9��9��9؇�9���9���9���9Z��9���9��9���9���9ѓ�9��9O��9��9���9�}�9t�9'q�9<m�9�h�97i�9�h�9�i�9x   x   \l�9o�9�r�9[t�9iy�9���96��9n��9H��9m��9Ȓ�9Ә�9���9u��9��9;��9֒�9H��9H��9^��9ӄ�9�9Qz�9t�9�q�9;p�9�l�9�j�9.k�9�j�9x   x   �s�9�o�9Xw�9�}�9���9���9.��91��9&��9~��9ϔ�9���9��9x��9���9���9a��9C��9��9V��9c��9���9�|�9�w�9�o�9�r�9Vq�9Up�9�o�9�q�9x   x   &{�9�x�9�~�9��95��9-��9Ɋ�9(��9��9���9M��9>��9���9��9���9��9���9ي�9
��9��9���9��9D�9Fy�9�z�9{�9�v�9@x�9(w�9Vz�9x   x   �{�9��9z��9��9n��91��9#��9ϓ�9��9ˑ�9ŗ�9J��9ٗ�9ї�9���9��9���9P��9d��9���9$��9���9�~�9�{�9\|�9�y�9u�9_�9�y�9�{�9x   x   c��9���9���9Շ�9I��9'��9��9!��9e��9/��9B��9œ�93��9��94��9ڒ�9}��9���9]��9χ�9N��9͋�9���9ڇ�94��9��9��9��9��9���9x   x   ��9=��9Ɛ�9���9n��9y��9���9ȑ�9)��9ݗ�9^��9���9���9���9���9Y��9���9��9e��9D��9���9���9���9��9I��9`��9f��9���9*��9ӏ�9x   x   ��9s��9͘�9���9˒�9˔�9N��9×�9?��9e��9	��9���9{��9!��9���9��9b��9��9��9��9��9ӓ�9"��9Q��9}��9���9N��9ܒ�9N��9��9x   x   ֗�9���9H��9���9Ԙ�9���9>��9H��9���9���9���9��9���9��9ך�9Ә�9���9Ж�9���9֖�9���9��9s��9���9H��9���9���9���9���9ו�9x   x   ���9���9���9[��9���9��9���9ۗ�93��9���9{��9 ��9���9V��9?��9���9Ě�9���9A��9!��9���9���9��9���9B��9w��9���9���9���9L��9x   x   1��9��9���9���9k��9v��9��9͗�9���9���9��9��9U��9ɛ�9q��9��9]��9���9P��9Ҥ�9���9���9ˤ�9���95��9`��9���9��9v��9̥�9x   x   ��9G��9���9��9��9���9���9���94��9���9���9Ԛ�9A��9r��9���9i��9Ȣ�9��9��98��9���9���9��9���9��9׮�9��9D��9���9m��9x   x   £�98��9?��9���9@��9���9��9��9֒�9^��9��9֘�9���9��9h��9ˢ�9���92��9���9ү�9���9���9���9	��9w��92��9_��9߮�9���95��9x   x   ���9���9���9���9ے�9]��9���9���9z��9~��9d��9���9Ú�9^��9̢�9���9���9-��9,��9���9���9���9���9���9?��9��9\��9@��9��9/��9x   x    ��9M��9R��9ӓ�9J��9C��9ي�9S��9���9��9��9ϖ�9���9���9���94��9-��9���9C��9���9y��9���9$��9���9?��9'��93��9T��9��9���9x   x   i��9w��9e��9��9J��9	��9��9^��9_��9g��9��9���9A��9N��9��9���9,��9G��9ֵ�9m��9̽�9;��9W��9���9a��9N��9��9���9���9��9x   x   ��9I��9F��9U��9_��9[��9���9���9ׇ�9J��9��9ߖ�9(��9Ѥ�9;��9ү�9���9���9h��9c��9���9u��9L��9��9��9���9v��9S��9��9���9x   x    ��9��9��9��9ք�9d��9���9#��9N��9���9��9���9���9���9���9���9���9���9̽�9���9���9��9F��9���9���9.��9H��9J��9��9˕�9x   x   ��9���9v��9���9Ā�9���9��9���9ы�9���9ؓ�9��9���9���9���9���9���9���93��9x��9��9\��9��9U��9���9���9���9���9���9ʓ�9x   x   Q��9V�9��9�}�9Tz�9�|�9F�9�~�9���9���9+��9x��9	��9Τ�9��9���9���9'��9R��9K��9@��9ܾ�9¶�9���9��9��9~��9���9|��9���9x   x   �|�9x�9w�9t�9t�9�w�9Fy�9�{�9��9��9V��9���9���9���9���9��9���9���9���9��9���9P��9���9���9_��9u��9��9O��9͉�9B��9x   x   Tz�9Hq�9�q�9+q�9�q�9�o�9�z�9_|�9:��9K��9���9O��9D��97��9��9|��9A��9C��9]��9��9���9���9��9c��9I��9���9H��9E��9M��9#|�9x   x   �r�9+o�9}m�9@m�9=p�9�r�9{�9�y�9��9`��9���9���9{��9d��9ٮ�95��9��9(��9I��9���9.��9���9��9v��9���9ю�9���9.��9By�9{�9x   x   �l�9mi�9d�9�h�9 m�9^q�9�v�9x�9��9e��9N��9���9���9���9��9d��9[��90��9���9|��9F��9���9y��9��9F��9~��9���9I�96w�9�q�9x   x   pi�9�d�98f�95i�9�j�9Vp�9Ex�9d�9��9���9��9���9���9��9G��9��9C��9W��9���9T��9L��9���9���9R��9I��93��9L�9�x�9�o�9Zj�9x   x   	d�9a�9}c�9�h�9-k�9�o�9'w�9�y�9��9*��9S��9���9���9y��9���9���9��9��9���9��9��9���9{��9ʉ�9H��9Dy�9/w�9�o�9/l�9 i�9x   x   �_�9�_�9;^�9�i�9�j�9�q�9Wz�9�{�9���9ԏ�9��9ܕ�9M��9Υ�9r��99��90��9���9��9���9Ε�9ȓ�9���9=��9|�9{�9�q�9Zj�9i�9\]�9x   x   1��9���9q��95��9J��9Y��9���9���9��9/��9���9A��9���9B��9���9���9���9���9��9��9���9<��9��9'��9g��9��9���9���9���9͡�9x   x   ���9��9T��9��9��9A��9���9���9���9���9`��9��9���9���9���9H��9���9.��9���9���9���9d��9[��9f��9��9���9��98��9%��9ۡ�9x   x   q��9U��9,��9&��9Q��9C��9f��9��9Q��9w��9��9���9 ��9)��9���90��9<��9��90��9���9���9��9p��9��9��9¯�9v��9~��9a��9��9x   x   /��9��9#��9G��9ؼ�9���9���9��9���9���9���9���9���9G��9<��9[��9v��9���9���9'��9M��9���9N��9���9���9z��9j��9ԥ�9���9Χ�9x   x   J��9��9K��9ڼ�9���9���9n��9���9���9��9/��9���9���91��9���94��9���9���90��95��9���9���9+��9˼�9��9���9��9���9��9��9x   x   X��9H��9C��9���9���9��9Z��9~��9���9���92��9X��9���9q��98��9���9��9���9���9h��9���9���9O��9v��9 ��9���9H��9��9 ��9��9x   x   ���9���9a��9���9k��9[��9>��9'��9R��9��9��9���9���9M��9��9t��9s��9���9x��9���9���9)��9?��9���9��9͸�9ϻ�9̳�9���94��9x   x   ���9���9��9��9���9��9(��9���9r��9���9X��9S��9���9���9���9���9G��9���9���9���9���9~��9��9*��9���9V��9*��9��9���9���9x   x   !��9���9K��9���9���9���9T��9p��9���9��9���9���9t��9���9���9X��9V��9:��9���9���9���9���9>��9���9R��9���9���9���9Q��9���9x   x   +��9���9u��9���9��9���9��9���9��9���9R��9A��9��9k��9:��9��9���9���9���9���9���9��9���9���9���9|��9���9��9���9���9x   x   ���9^��9��9���9.��93��9��9]��9���9W��9%��9q��9/��9��9���9���9_��95��9n��9��9Q��9���9K��9���9i��9���9���92��9���9���9x   x   <��9��9���9���9���9S��9���9T��9��9G��9x��9���9���9/��9��9���9���9W��9���9���9���9���9{��96��9���9.��9���9 ��9���9G��9x   x   ���9���9���9���9���9���9���9���9r��9��9,��9���9��9���9+��9���9��9���9���9���9W��94��96��95��9=��9p��9\��9P��9-��9���9x   x   >��9���9%��9C��93��9u��9M��9���9���9k��9��93��9���9���9���9z��9���9>��9���9U��9���9)��9���9���9���9���9���9���9��9���9x   x   ���9���9���9=��9���93��9��9���9���9:��9���9��9*��9���9|��9���9H��9��9��9U��9��9��9N�9���9� �9#�9���9:��9���9p��9x   x   ���9C��9+��9[��93��9���9s��9���9Y��9��9���9���9���9{��9���9���9���9���9p��9S��9$ �9?�9��9��9��9' �9���9���9D��9���9x   x   ���9���98��9n��9���9��9z��9E��9\��9��9a��9���9��9���9F��9���9B��9� �9�9D�9I
�9��91�9%�9�
�9��9��9! �9}��9���9x   x   ���92��9	��9���9���9���9���9���9B��9���9>��9^��9���9B��9	��9���9� �9��9�	�9W�9��9��9%�9a�9��9	�9�9� �9���9���9x   x   ��9���95��9���9.��9���9t��9���9���9���9r��9���9���9���9��9r��9�9�	�9��9��9��9��9�9!�9��9;	�9�9c��9���9���9x   x   ��9���9���9*��99��9j��9���9���9 ��9���9 ��9���9���9W��9W��9R��9G�9S�9��9X�9��9��9,�96�9(�9��9���97��98��9���9x   x   ���9���9���9O��9���9���9���9���9���9���9T��9���9X��9���9��9( �9J
�9��9��9��9��92�9��9&�9g
�9���9���9���9���9��9x   x   <��9e��9��9���9���9���91��9���9���9	��9���9���98��9,��9��9A�9��9��9��9��91�9��9�9��9��9��9	��9���9���9���9x   x   ��9^��9r��9N��9*��9K��9F��9��9@��9���9M��9���97��9���9K�9��95�9$�9&�9+�9��9�9T�9L�9h�9+��9C��9>��9���9&��9x   x   )��9j��9��9���9̼�9w��9���9(��9���9���9���98��96��9���9���9��9%�9b�9�96�9'�9��9P�9���90��9c��9���9Y��9���9��9x   x   j��9��9��9���9��9!��9��9���9T��9���9l��9���9@��9���9� �9��9�
�9��9��9-�9c
�9��9f�9+��9'��9���9��9���9���9���9x   x   ��9��9���9z��9���9���9ٸ�9\��9���9���9���96��9u��9���9#�9. �9��9	�9A	�9��9���9��9-��9d��9���9���9��9A��9���9a��9x   x   ���9��9|��9j��9��9G��9л�9,��9���9���9���9���9a��9���9���9���9��9�9�9 �9���9��9D��9���9��9��9l��9}��9���9~��9x   x   ���98��9��9ԥ�9���9��9ʳ�9��9���9��97��9%��9Q��9���9;��9���9! �9� �9_��96��9���9���9;��9Y��9���9>��9}��9/��9k��9���9x   x   ���9 ��9b��9���9��9)��9���9���9X��9���9���9���9-��9��9���9D��9��9���9���9?��9���9���9���9���9���9���9���9o��9ެ�9��9x   x   ס�9ߡ�9���9ͧ�9��9��9:��9���9���9���9���9D��9���9���9m��9���9���9���9���9���9��9���9&��9 ��9���9_��9���9���9��9e��9x   x   !��9���9���9��9���9���96��9;�9��9��9*�9�/�9�;�98>�9�<�9HE�9�<�9)>�9�;�9>1�9�*�9��9��9F
�9���9��9N��9��9���9.��9x   x   ���9%��9���9���9l��9���9�9�9��9�#�9�*�9�1�9�8�9�;�9
=�9C>�9�:�9#9�9�1�9>)�9d"�9��9��9��9���9��9��9j��9���9��9x   x   ���9���9E��91��9��96��9f�9��9w�9�#�9�+�9�0�903�9�;�9z8�9�:�9�3�9T0�9d,�9!&�9��9��9�	�9T��9 ��9���9���9��9&��9O��9x   x    ��9���93��9
��9���9^�9��9��9; �9�'�9�-�9�/�9�4�9[6�9+6�9}5�9�.�9y.�9&�9b�9C�9��9S�9 ��9!��9���9$��9F��9���9f��9x   x   ���9e��9��9���9�9,
�9��9��9��9�#�9�)�9Q/�9�3�9`3�9�3�9/�9w*�9�#�9!�9/�9��9�	�9�9���9���9���9���9���9���9}��9x   x   ���9���92��9Z�9+
�9P�9��9)!�9t#�9�&�9�(�9X/�9N3�9k3�9�.�9)�9�%�9�"�9V �9��9��9T�9��94��9���9���9���9���9���9���9x   x   0��9�9i�9��9��9��9��9��9�%�9�,�9e+�9Z.�9+�9�.�9�+�9U,�9x'�9"�9��9��9��9t�90
�9��9W��9��9b��9���9>��9���9x   x   6�9�9��9��9��9(!�9��9�"�9z*�9e+�9(-�9,�9�+�9�,�9�+�9�)�9B"�9s�9�!�9[�9��9#�9��9��9�	�9�	�9��9w
�9Z
�9r
�9x   x   ��9��9s�99 �9��9w#�9�%�9x*�9�%�9�(�9�0�9;2�9m1�9�(�9�&�9�*�9�%�9�!�9Z �9� �9�9��9E�91�9B�9��9$�9��9��9M�9x   x   ��9�#�9�#�9�'�9�#�9�&�9�,�9a+�9�(�9.0�9Y.�9�-�90�9�'�91+�9,�9�'�9�#�9�$�9�%�9�"�9i�9��9�9�96�9J�9R�9��9F�9x   x   
*�9�*�9�+�9�-�9�)�9�(�9c+�9$-�9�0�9U.�9�%�9W.�9�1�9P-�9�+�9�'�9=)�90�9�,�9�)�9+�9�(�9�.�9�(�9�'�9�'�9�'�9�(�9.�9�(�9x   x   �/�9�1�9�0�9�/�9L/�9U/�9Y.�9",�9=2�9�-�9W.�9n1�9�+�9�-�9Z0�9�0�9�-�9�/�9i1�9�0�971�9�.�9�0�9�3�9 5�9�4�9{4�9C/�9�/�9�2�9x   x   �;�9�8�933�9�4�9�3�9J3�9+�9�+�9r1�90�9�1�9�+�9�+�9�2�9�1�9R6�9�4�99�9<�9�:�9^?�95;�9�<�9?�91;�9�>�9k=�9�<�9{<�9�;�9x   x   7>�9�;�9�;�9\6�9]3�9l3�9�.�9�,�9�(�9�'�9T-�9�-�9�2�9�5�9�5�9:�9;�9�=�9�B�9�A�9�G�9�G�9I�9mJ�9�J�9�H�9vF�9�H�9�B�9�B�9x   x   �<�9
=�98�9.6�9�3�9�.�9�+�9�+�9�&�9.+�9�+�9b0�9�1�9�5�9�9�9�=�9�=�96C�9�J�9[K�9aP�9KO�9.Q�9�U�9&Q�9�P�9'O�9rL�9�I�9C�9x   x   FE�9A>�9�:�9|5�9/�9)�9R,�9�)�9�*�9�,�9�'�9�0�9U6�9:�9�=�9�C�9�H�9&I�9�P�9�W�9�[�9;]�9K_�9h_�9�[�9�\�9�W�9P�9�J�9I�9x   x   �<�9 ;�9�3�9�.�9{*�9�%�9v'�9B"�9�%�9(�9C)�9�-�9�4�9;�9�=�9�H�9>R�9�U�9'Z�9�Y�9^�9pc�9ha�9)e�9�]�9�Z�9�Z�9�U�9IP�9�G�9x   x   $>�99�9T0�9w.�9�#�9�"�9!�9t�9�!�9�#�90�9�/�99�9�=�9;C�9)I�9�U�9�\�99_�9nb�9�e�9�i�9%g�9�e�9�a�9�^�9j\�9oU�9L�9�C�9x   x   �;�9�1�9c,�9&�9!�9W �9��9�!�9\ �9�$�9�,�9k1�9
<�9�B�9�J�9�P�9(Z�98_�9�j�96k�9
i�9{p�9aj�9Yk�9�k�9�_�9TZ�9�O�9lH�9�B�9x   x   >1�9B)�9 &�9_�9/�9��9��9]�9� �9�%�9�)�9�0�9�:�9�A�9^K�9�W�9�Y�9sb�96k�9�l�9�n�9o�9k�9�j�9�a�9�Y�9�X�9=L�9�C�9q:�9x   x   �*�9j"�9��9D�9��9��9��9��9�9�"�9+�9:1�9f?�9�G�9dP�9�[�9^�9�e�9i�9�n�9^k�9�n�9k�9�e�9U_�9�Z�9�O�9VG�9b=�9�1�9x   x   ��9��9��9��9�	�9[�9u�9'�9��9p�9�(�9�.�9<;�9�G�9RO�9B]�9rc�9�i�9�p�9o�9�n�9�o�9�g�9c�9*]�9�P�9�G�9<�9#0�9<(�9x   x   ��9��9�	�9R�9!�9��90
�9��9I�9��9�.�9�0�9�<�9I�9.Q�9P_�9na�9'g�9bj�9k�9k�9�g�9�c�9n^�9�P�9H�9�<�9�/�9�-�9K�9x   x   I
�9��9Z��9"��9���9<��9��9��9=�9�9�(�9�3�9?�9vJ�9�U�9e_�9.e�9�e�9[k�9�j�9�e�9c�9m^�9~W�9J�9@�9�3�9B)�9�9��9x   x   ���9���9��9!��9���9���9]��9�	�9E�9�9�'�95�9/;�9�J�9+Q�9�[�9�]�9�a�9�k�9�a�9Z_�9(]�9�P�9J�9 ;�9�4�9�(�9��9��9|�9x   x   ��9��9���9���9���9���9��9�	�9��9;�9�'�9�4�9�>�9�H�9�P�9�\�9�Z�9�^�9�_�9�Y�9�Z�9�P�9}H�9@�9�4�9�'�9)�9n�9g	�9#��9x   x   M��9��9���9!��9���9���9e��9��9#�9R�9�'�94�9o=�9�F�9/O�9�W�9�Z�9m\�9VZ�9�X�9�O�9�G�9�<�9�3�9�(�9+�9��9�
�9���9���9x   x   ��9r��9��9K��9���9���9���9}
�9��9S�9�(�9C/�9�<�9�H�9wL�9P�9�U�9qU�9�O�9@L�9YG�9<�9�/�98)�9��9n�9�
�9"��9���9���9x   x   ���9���9(��9���9���9���9A��9`
�9��9��9.�9�/�9�<�9�B�9�I�9�J�9GP�9	L�9nH�9�C�9b=�9$0�9�-�9�9��9d	�9���9���9���9��9x   x   4��9��9M��9k��9y��9���9���9t
�9U�9S�9�(�9�2�9�;�9�B�9C�9I�9�G�9�C�9�B�9u:�9�1�98(�9O�9��9}�9��9���9|��9��9K��9x   x   �!�9b�9��9�)�9�+�9�:�9F�9�Q�9�a�9ck�9Jq�9�9���9&��9���9x��9��9��9X��9Հ�9�p�9Nk�9a�9�O�9�F�9'<�9�+�9p(�9� �9��9x   x   ]�9��9}#�9�*�93�9�;�9�B�9�P�9�]�98m�9�y�9W��9��9b��9ώ�9��9���9��9��9Sy�9Hm�9K]�9�S�9�B�9:�9�2�9�+�9�"�9��9e�9x   x   ��9w#�99)�92�9�;�9�C�9�Q�9Z�9�c�9�j�9�w�9|�9ւ�9F��9���9���9߃�9i|�9Sw�9�k�9�d�9%X�9�O�9�D�9�<�9=1�9�)�9�$�9��9��9x   x   �)�9�*�92�9/7�9�=�9-M�9�S�9g_�9�d�9ho�9z�9~�9<��9x��9��9S��9{|�9{�9So�9$b�9Qa�9�T�9gM�9;<�9�7�9�1�9�)�9�)�9%�9&�9x   x   �+�93�9�;�9�=�9�N�9�S�9�X�9�c�9'j�9t�9oz�9��9��9W��9��9*��9�z�9�r�9�l�9�c�9qV�9T�9ZO�9/=�9�;�94�9=+�9�)�97+�9�(�9x   x   �:�9�;�9�C�9(M�9�S�9pX�9D`�9�n�9�q�9�v�9%}�9�~�9y�9iy�9�}�9,}�9w�9�p�9�m�9�a�9�Y�9R�93N�9�C�9Z:�9l;�9�3�9�2�9�3�9�4�9x   x   F�9�B�9�Q�9S�9�X�9H`�9�e�9�p�9�r�9�u�9{�9���9={�9}��9�{�9~t�9:t�9�p�9�e�9/_�9}Y�9FT�9�O�9�C�9�E�9~C�9�;�9�>�9G;�9C�9x   x   �Q�9�P�9Z�9d_�9�c�9�n�9�p�9�t�9w�96x�9O~�9�}�9�}�9~�9�x�9xv�9�s�9r�9�n�9�c�9�^�9�Z�9%Q�9�Q�9fN�9�E�9�J�9fJ�9!F�9�N�9x   x   �a�9�]�9�c�9�d�9(j�9�q�9�r�9w�9�{�9�|�9�x�9�v�9y�9�{�9C|�9�w�9�r�9Rp�9�k�9�d�9c�9Y^�9�`�9S[�9	Y�9�W�9<V�9�X�9EX�9OZ�9x   x   \k�97m�9�j�9do�9t�9�v�9�u�98x�9�|�9�z�93|�9B{�9|�9�|�9=w�9v�9�w�9�s�9�l�9ol�9�l�9Wk�9�j�9�b�9�j�9wh�9�g�9�i�9d�9j�9x   x   Aq�9�y�9�w�9z�9jz�9$}�9{�9H~�9�x�96|�9Հ�9|�9�w�9�9�{�9�{�9[z�9�{�9Fx�9-x�9�q�9Ut�9uv�9�q�9�u�9�r�9�v�9�q�94v�9�s�9x   x   �9U��9|�9�}�9��9�~�9���9�}�9�v�9C{�9|�9�v�9�}�9���9w�9��9�{�9e{�9���9���9R�9ǃ�9j��9O��9���9��96��9H��9ل�9k��9x   x   ���9��9΂�9:��9��9y�9?{�9�}�9!y�9|�9�w�9�}�9h{�9ey�9�}�9_��9���9ȃ�95��9��9��9���9i��9��9َ�9��9���9C��9���9܋�9x   x    ��9]��9=��9v��9T��9ky�9}��9~�9�{�9�|�9�9���9dy�9���9a��9ǈ�9���9Ǝ�9���9v��9ԗ�9���9ߛ�9��9ʟ�9Ú�9���9��9��9>��9x   x   ���9ˎ�9���9��9��9�}�9�{�9 y�9D|�9?w�9�{�9t�9�}�9_��9v��9e��96��9Ɨ�99��9ܞ�9���9��9e��9���9���9|��9��9Y��9}��9Z��9x   x   t��9��9���9T��9)��9)}�9�t�9v�9�w�9v�9�{�9��9c��9Ɉ�9m��9��98��9���9p��9«�9s��9t��9>��9���9`��9ȳ�9���9���9��9̝�9x   x   ��9���9ރ�9||�9�z�9w�97t�9�s�9�r�9�w�9\z�9�{�9���9���97��97��9��9R��9W��9���9ۻ�9��9 ��9P��9e��9Q��9���9~��9s��9��9x   x   ��9��9h|�9�z�9�r�9�p�9�p�9r�9Qp�9�s�9�{�9f{�9̓�9ʎ�9�9���9W��9��9T��9��9���9���9@��9���9���9��9ծ�9��9%��9=��9x   x   Y��9��9Ow�9Zo�9�l�9�m�9�e�9�n�9�k�9�l�9Ix�9���96��9���9=��9m��9Y��9Q��94��9:��9V��9���9���9��9V��9h��9���99��96��9S��9x   x   ڀ�9Vy�9�k�9&b�9�c�9�a�90_�9�c�9�d�9sl�93x�9���9��9x��9��9ǫ�9���9"��96��9i��9U��9���9���9���9ϼ�9��9���9���9��9̊�9x   x   �p�9Gm�9�d�9Qa�9uV�9�Y�9�Y�9�^�9c�9�l�9�q�9W�9��9՗�9���9p��9ػ�9���9T��9V��9���9p��9���9��9���9��9"��9���9}��9]�9x   x   Lk�9K]�9)X�9�T�9T�9R�9GT�9�Z�9^^�9]k�9Wt�9Ƀ�9���9���9��9z��9��9���9���9���9o��9���9���9���9��9ԥ�9h��9���9U��9u�9x   x   a�9�S�9�O�9hM�9_O�9:N�9�O�9/Q�9�`�9�j�9|v�9l��9n��9���9g��9A��9&��9A��9���9���9���9���9���9���96��9��9ב�9���9t�9k�9x   x   �O�9�B�9�D�9?<�93=�9�C�9�C�9�Q�9T[�9�b�9�q�9X��9��9��9���9���9T��9���9��9���9��9���9���9���9%��9ޑ�9���9Ms�9$d�9�Z�9x   x   �F�9:�9�<�9�7�9�;�9Z:�9�E�9kN�9Y�9�j�9�u�9���9ݎ�9Ο�9���9g��9h��9��9[��9Ҽ�9Ľ�9��9>��9,��9���9��9hu�9�i�9�W�9tP�9x   x   ,<�9�2�9G1�9�1�9 4�9r;�9�C�9�E�9�W�9�h�9�r�9��9���9�9��9ȳ�9V��9��9j��9��9��9֥�9��9ޑ�9��9{t�9�g�9�Y�93E�9�A�9x   x   �+�9�+�9�)�9�)�9?+�9�3�9�;�9�J�9CV�9�g�9�v�9=��9���9���9��9���9���9׮�9��9���9"��9f��9Ց�9���9fu�9�g�93V�9%J�9b=�9�3�9x   x   s(�9�"�9�$�9�)�9�)�9�2�9�>�9nJ�9�X�9�i�9�q�9O��9B��9��9_��9���9���9��98��9���9���9���9���9Ps�9�i�9�Y�9%J�9�=�9�2�9�)�9x   x   � �9��9��9%�96+�9�3�9K;�9(F�9JX�9�d�97v�9��9���9��9~��9��9z��9'��94��9��9}��9W��9t�9'd�9�W�97E�9a=�9�2�9%+�9�%�9x   x   ��9b�9��9
&�9�(�9�4�9C�9�N�9LZ�9j�9�s�9q��9ߋ�9?��9]��9͝�9"��9B��9U��9Ί�9_�9u�9 k�9�Z�9tP�9�A�9�3�9�)�9�%�9G�9x   x   M�9U�9xY�9k`�9�k�9wt�9	��95��9z��9ķ�9
��9���96��9z��9���9���9���9��9I��9���9m��9���9���9���9��9+v�9�j�9z_�9%[�98U�9x   x   
U�9z`�9*\�99j�9Ds�9�~�9���9<��9���9���9���9��9)��9���9���9���9���91��9���9���9J��9V��9���9��9/}�9�s�9k�9"\�9�^�9�T�9x   x   |Y�9$\�90`�9�m�9�w�9��9���9���9(��9���9���9���9o��9���9���9���9Q��9/��9���9���9'��9+��9��9���9�v�9�l�9`�9�\�9�Z�9iX�9x   x   l`�95j�9�m�9�t�9σ�9ш�9͗�9ͨ�9���9���9��9���9m��9���9���9���9���9���9.��9ʵ�9Ū�9h��9p��9���9�u�9n�9�i�9�_�92_�9�`�9x   x   �k�9Bs�9xw�9҃�9���9Γ�9p��9��9ŷ�9��91��9���9V��9C��9���9���9���9���9��9%��9W��9���9��9$��9Pv�9�s�9dl�9rg�9g�9�f�9x   x   wt�9�~�9���9ш�9ԓ�9���9���9���93��9���9���9f��9W��9#��9{��9���9���9��9*��9o��92��9�9u��9ǈ�9�~�9Zt�9�u�9�u�9�u�9�v�9x   x   ��9���9���9ȗ�9k��9���9���9��9���9'��9Q��9I��9���9���9���9���9��9}��9Գ�9���9$��9"��9���9���9Ĉ�9���9���9�9���9x��9x   x   .��96��9���9Ψ�9��9���9��9}��9���9���9���9���9���9���95��9��9���9���9���9���9]��9y��9���9���9(��9���9��9=��9P��9ϐ�9x   x   v��9���9 ��9���9���91��9���9���9���9���9���9v��9���9W��9���9~��9���9���9���9���9L��9��9j��9���9���9��9���9��9���9&��9x   x   ���9���9���9���9��9���9#��9���9���9'��9-��9���96��9��9���9v��9w��9���9Z��9���9���9��9)��9��9F��9-��9ư�9���9��9���9x   x   ��9���9���9��94��9���9N��9���9���9/��9|��9���9���9��9���9��9:��9���9Z��9Z��9���9h��9
��9���9���9���9$��9��9���9��9x   x   |��9��9���9���9���9Z��9B��9���9t��9���9���9��9���9h��9w��9$��9��9���9���9=��9J��9j��9���9;��9+��9���9���9��9C��9F��9x   x   3��9)��9p��9o��9W��9O��9���9���9���94��9���9���9���9���9!��9���9���9���9���9��9���9���9���9���9~��9���9#��9��9;��9���9x   x   v��9���9���9���9E��9!��9���9���9X��9��9��9q��9���9��9���9���9!��9���9H��9S��9(��9���9I��9��9���9��9���9��9J��9���9x   x   ���9���9���9���9���9s��9���92��9���9���9���9}��9%��9���9���9���9���9���90��9h��9P��90�9�9���9��9c�9���9���9���9���9x   x   ���9���9���9���9���9���9���9��9��9y��9��9'��9���9���9���9y��9,��9���9j�9��9&�9��9��9��9��9��9��9P�9���9���9x   x   ���9���9M��9}��9���9���9��9���9���9y��9;��9��9���9!��9���9+��9��9.�9��9�94�9�9c!�9O�9Z�97�9��9��9���9���9x   x   ��95��95��9���9���9��9���9���9���9���9���9���9���9���9���9���92�9r�9��9��92�9�#�9E#�9�9��9��9��9��9���9���9x   x   I��9���9���9+��9���9-��9г�9���9���9[��9`��9���9���9N��96��9k�9��9��9/�9�$�9�)�9�+�9*�92$�9��9��9Q�9� �9!��9v��9x   x   ���9���9���9ε�9'��9r��9���9���9���9���9Z��9A��9 ��9W��9i��9��9�9��9�$�9 0�9J+�9�*�950�9�%�9�9v�9��9���9?��9���9x   x   n��9N��9(��9ʪ�9X��95��9+��9b��9U��9���9���9O��9���9.��9R��9-�9:�97�9�)�9L+�9�%�9C+�9�(�9�9 �9��9���9���9��9���9x   x   ���9Z��9-��9o��9��9ǒ�9,��9}��9��9!��9s��9o��9���9���93�9��9�9�#�9�+�9�*�9>+�9�,�9D#�9�9��9��9���9j��9���9���9x   x   ���9���9���9s��9���9x��9���9���9o��93��9��9���9���9R��9%�9��9j!�9J#�9$*�990�9�(�9I#�9#�9o�9t�93��9���9	��9���9ز�9x   x   ���9��9���9���9'��9ˈ�9���9���9���9��9���9:��9���9(��9��9��9S�9#�92$�9�%�9�9�9q�9���9���99��9���9���9m��9/��9x   x   ��99}�9�v�9�u�9Zv�9�~�9Έ�92��9���9Q��9���9.��9���9���9��9��9X�9��9��9�9��9��9l�9���9���9C��9���9���9��9���9x   x   .v�9�s�9�l�9n�9�s�9\t�9���9���9���93��9���9���9���9��9f�9��9=�9��9��9u�9��9��90��9;��9G��9��9Y��9Y��9���9=��9x   x   �j�9k�9`�9�i�9gl�9�u�9���9��9���9ǰ�9+��9���9.��9���9���9��9��9��9R�9��9���9��9���9���9���9S��9?��9Վ�9Έ�9*u�9x   x   _�9!\�9�\�9�_�9xg�9�u�9�9A��9��9���9��9��9��9��9���9R�9��9��9� �9���9���9k��9��9���9���9S��9Ԏ�9�|�9�u�9�h�9x   x   *[�9�^�9�Z�98_�9g�9�u�9���9Q��9���9��9���9K��9@��9U��9���9���9���9���9'��9F��9��9���9���9m��9��9���9ʈ�9�u�9Rf�9�_�9x   x   =U�9U�9gX�9�`�9�f�9�v�9z��9֐�91��9��9��9J��9���9���9���9���9���9���9y��9���9���9���9ղ�93��9���9;��9+u�9�h�9�_�9�W�9x   x   F��9;��9��9W��9���9���9��9���9��9� �9p�9F!�9�4�9~7�9�=�9�C�9�?�9�8�9!3�9�!�9~�9���9���9���9���9���9���9ƙ�9���9B��9x   x   8��9���9=��9E��9���9W��9C��9���9'��99�9��9"�9\+�9U1�9�:�99�9d/�9�+�9�"�9��9�9 ��9���9���9��9ɰ�9��9ޘ�9�9Ƌ�9x   x   ��9>��9v��9��9��9i��9&��9S��9��9�	�9d�9( �9�$�9i.�95�91�9%�9��9��9	�9���9���9���9��9��9Z��9���95��9���9֒�9x   x   P��9G��9��9���9m��9.��9M��9E��9���9I
�9��9� �9p)�9�'�9b&�9X(�9s �9��91�9��9���9���9��9���9���9��9���9˙�9R��9Y��9x   x   ���9���9��9l��9���9��9g��9���9v�9��9u�9f!�9�$�9��9+%�9�"�9��9��9B�9��9���9m��9Q��9���9˵�9>��9��9e��9l��9��9x   x   ��9X��9k��9+��9��9��9i��9T�9��9��9*�9#�9��9��9@"�9p�9��9�9�9���9!��9���9>��9_��9��9��9���9��9`��9��9x   x   ��9?��9%��9K��9d��9g��9�9-�9��9R�9��9��9��9.�9� �9�9?�9��9; �9���9���9H��9��9���9���9���9ɽ�9���9��9��9x   x   ���9���9T��9E��9���9U�9,�9��9��9��9��9��9�9�9��9��9��9��93�9p��9C��9��9���9l��9���9���9���99��9;��9!��9x   x   ��9#��9��9���9v�9��9��9��9��9��9�!�9��9�!�9:�9��9��9��9��9��9���9@��9���9��9���9���9G��9Y��9���9���9���9x   x   � �94�9�	�9E
�9��9��9W�9��9��9��9h�9�9��9��9{�9�9>�9G�9L
�9�
�9��9U �9���9� �9���9}��9<��9���9���9���9x   x   j�9��9[�9��9p�9(�9��9��9�!�9c�9,�9!�9d�9�9 �9��96�9��9<�9 �9��9��9Y�9L�9��9��9��9��9��9��9x   x   A!�9"�9% �9� �9g!�9#�9��9��9��9�9!�9 �9��9��9_"�9�"�9  �9 �9g#�9�!�9!�9m%�9g&�9S(�9'�9�%�9�'�9�'�9�$�9 �9x   x   �4�9V+�9�$�9i)�9�$�9��9��9��9�!�9��9f�9��9'�9! �9�$�9�(�9c%�9+�9�3�9�4�9�3�9N<�9�;�9:�9�;�9`;�9G;�9�:�9�5�9e5�9x   x   {7�9J1�9d.�9�'�9��9��9-�9}�9<�9��9�9��9 �9��9�'�9N/�9�0�9�7�9�A�9TG�9�F�9[I�9�L�90O�9O�9L�9NJ�9�G�9�E�90@�9x   x   �=�9�:�95�9]&�9(%�9A"�9� �9��9��9�9 �9^"�9�$�9�'�9�4�9�9�9�>�9�E�9�I�9�S�9O[�9
Y�9�_�9c�9�_�9�Y�9�Z�9�R�9�L�9�F�9x   x   �C�99�91�9V(�9�"�9s�9��9��9��9�9��9�"�9�(�9U/�9�9�9OD�9wP�9?Y�9�Z�9�f�9+n�9}o�9Uo�9�o�9�o�9!m�9fh�9�Z�9IV�9Q�9x   x   �?�9_/�9%�9o �9��9��9>�9��9��9>�9<�9 �9j%�9�0�9�>�9�P�9�Y�9�b�9�k�9ur�9��9���9+~�9 ��9T��9jr�9�j�9uc�9_[�9sP�9x   x   �8�9�+�9��9��9�9�9��9��9��9K�9��9 �9+�9�7�9�E�9?Y�9�b�9�j�9�r�9���9C��9���9$��9��9΁�9�r�9�j�9vb�9zW�9�D�9x   x    3�9�"�9��91�9D�9�9B �99�9��9Q
�9C�9q#�9�3�9�A�9�I�9�Z�9�k�9�r�9��9'��9���9�9Í�9���9R��9�s�9sj�9�Z�9�L�9�@�9x   x   �!�9��9	�9��9��9��9��9v��9���9�
�9�9�!�9�4�9TG�9�S�9�f�9rr�9���9'��9���9L��9���9<��9���9J��9Dr�9�h�9�Q�9F�9�5�9x   x   ��9�9���9���9���9"��9���9H��9K��9��9��9!�9�3�9�F�9W[�90n�9��9I��9���9F��9>��9%��9���98��9��9�l�9N[�9�G�9�4�9A �9x   x   ���9"��9���9���9q��9���9L��9��9���9X �9��9o%�9P<�9^I�9Y�9�o�9���9���9���9���9%��9���9ȇ�9��9�o�9BY�9�I�9�;�9�$�9��9x   x   ���9���9���9 ��9T��9F��9���9���9���9���9X�9o&�9�;�9�L�9�_�9Yo�91~�9$��9ō�9>��9���9Ç�9D�9�o�99`�9L�9;�9B'�9��95 �9x   x   ���9���9��9���9���9^��9���9t��9���9� �9U�9`(�9":�99O�9
c�9�o�9��9��9���9���98��9��9�o�9�a�9�O�9M;�9r(�9�9���9���9x   x   ���9���9��9���9ҵ�9��9���9���9���9���9��9'�9�;�9
O�9�_�9�o�9W��9ց�9Y��9P��9���9�o�9<`�9�O�9�:�9X&�93�9{��99��9V��9x   x   ���9ʰ�9_��9��9?��9��9���9���9H��9���9��9�%�9k;�9"L�9�Y�9.m�9nr�9�r�9�s�9Ir�9�l�9CY�9L�9N;�9Z&�9��9���9���9���9?��9x   x   ��9��9���9���9���9���9Ͻ�9���9e��9E��9��9�'�9J;�9TJ�9�Z�9kh�9�j�9�j�9sj�9�h�9K[�9�I�9;�9k(�96�9���9���9���9=��9��9x   x   ���9���91��9͙�9k��9��9���9B��9���9���9��9�'�9�:�9�G�9�R�9�Z�9{c�9~b�9�Z�9�Q�9�G�9�;�9D'�9�9|��9���9���9���9���93��9x   x   ���9ǎ�9���9X��9m��9d��9��9C��9���9���9��9�$�9�5�9�E�9�L�9OV�9`[�9W�9�L�9F�9�4�9�$�9��9���9=��9���9?��9���9$��9���9x   x   <��9Ë�9ג�9^��9��9��9��9!��9���9 �9��9 �9m5�90@�9�F�9Q�9vP�9�D�9�@�9�5�9A �9��94 �9���9T��9>��9��9.��9���93��9x   x   ���9���9G��9��9���9"��9�9D$�9L9�9Q�9;h�9�x�9��9_��9���9a��9���9��9c��9:x�9�h�9�P�9�9�9
$�9>�9;��9���9a��9���9���9x   x   ���9��9���9���9��9��9F�9�&�9�<�9 T�9gh�9:t�9a��9���9W��9Ԑ�9@��9g��9�u�9�g�9_T�9�<�9M&�9��9���9r��9h��9���9��9վ�9x   x   B��9���9R��9���9���9�	�9��90�9�G�9DW�9�i�9ct�9���9ԇ�9��9���9���9_s�9ci�9W�9�G�970�9�9�
�9��9x��9W��9J��9z��9��9x   x   ~��9���9���9���95��9o�9,$�9�;�9�N�9�U�9�m�9�p�9;}�9��9*��9T|�9�q�9�m�9�V�9�N�9�;�9�$�9o�9���9+��9,��9���9���9���9 ��9x   x   ���9��9���92��9��9��9/�9�G�9�P�9�]�9Gp�9�m�9�x�9�~�9�x�9Un�9�o�9]�95P�9�G�97.�9b�9��9	��9B��9���9��9��9���9���9x   x   !��9��9�	�9j�9��9i.�94>�9#L�9X�9�`�9l�9�o�9:s�9�s�9�o�9�j�9b�9lX�9cL�9?�9�-�9��9l�9
�9/��9S��96��9	��9���9��9x   x   	�9=�9��9$$�9/�97>�9�E�9�S�9�^�9�a�9�h�9s�9�v�9�q�97j�9vb�9]�9�S�9D�9�>�9/�9�#�9��9��9�
�9�9��9*�93��9��9x   x   =$�9�&�90�9�;�9�G�9L�9�S�9�X�9�d�9"h�95l�9�q�9s�9�l�9�f�9�d�9�Y�9*T�9jL�9OG�9$<�9"0�9'�9�$�9#�9��93�9��9��9%�9x   x   C9�9�<�9�G�9�N�9�P�9X�9�^�9�d�9�l�9tm�9yn�9|i�9�m�96m�9tm�9e�9�\�9�X�9hP�9�N�9�G�9><�9�8�9�3�9U0�9�0�96)�9�0�9�/�9%4�9x   x   Q�9T�9EW�9�U�9�]�9�`�9�a�9$h�9vm�9Ol�9zo�9Zo�9Om�9�m�9zf�9c�9�a�9�\�9�V�9W�9�T�9�Q�9M�9�F�9FK�9eH�9sG�9�K�9G�9�L�9x   x   ,h�9bh�9�i�9�m�9Cp�9l�9�h�92l�9}n�9}o�9-|�9Zo�9�l�9�l�9si�9<k�9�o�9n�9�h�9:h�9g�9�e�9�a�9/`�9�b�9k_�93c�9p_�9,a�9f�9x   x   �x�9;t�9bt�9�p�9�m�9�o�9s�9�q�9�i�9_o�9Zo�9�j�9xr�9�r�9�n�9�n�9iq�9�s�9�u�9=y�9z�9�|�9Qs�92z�9�y�9�y�9�y�9�t�9}�9!y�9x   x   ��9Z��9���98}�9�x�96s�9�v�9s�9�m�9Nm�9�l�9wr�9v�9$t�9ty�9�{�9���9���9��9���9���94��9���9��9ޒ�9���9���9�9���9܉�9x   x   ]��9���9Ӈ�9��9�~�9�s�9�q�9�l�98m�9�m�9�l�9�r�9't�91}�9��9Ĉ�9���9Ŕ�9Қ�9���9Ƣ�9F��9
��9ϭ�9V��9ݭ�9٫�9_��9K��9M��9x   x   ���9Q��9��9*��9�x�9�o�94j�9�f�9qm�9zf�9zi�9�n�9yy�9���9��9\��9)��9���9��9���9���9T��9���9���9C��9���9��9y��9ٳ�9��9x   x   _��9ΐ�9���9P|�9Rn�9�j�9zb�9�d�9�d�9c�9<k�9�n�9�{�9���9[��9���9��9���9���9���9��9���9w��9���9���9���9���9G��9N��9@��9x   x   ���9=��9���9�q�9�o�9b�9]�9�Y�9�\�9�a�9�o�9oq�9���9���9+��9��9��9&��9?��9���9���9��9���9��9��9���9g��99��9ױ�9C��9x   x   ��9e��9_s�9�m�9]�9nX�9 T�93T�9�X�9�\�9n�9�s�9���9ʔ�9���9���9%��9���9��9���9���9���9*��9���9���9���9���97��9T��9b��9x   x   d��9�u�9di�9�V�98P�9cL�9D�9pL�9oP�9�V�9�h�9�u�9 ��9ޚ�9��9���9C��9��9\��9��9
��9,��9/��9���9%��9f��9���9���9x��9���9x   x   8x�9�g�9W�9�N�9�G�9?�9�>�9UG�9�N�9W�9>h�9?y�9���9���9���9���9���9���9��9���9� �9F �9���9���9���9���9d��9���9���9���9x   x   �h�9_T�9�G�9�;�9C.�9�-�9'/�91<�9�G�9�T�9	g�9!z�9�9Ϣ�9���9��9���9���9	��9� �9L�9_ �9��9o��9+��9���9Ӽ�9*��9���9qy�9x   x   �P�9�<�9<0�9�$�9d�9��9�#�9+0�9J<�9�Q�9�e�9�|�9>��9O��9]��9���9��9���98��9N �9d �9q��9���98��9���9���9��9a��9�|�9�e�9x   x   �9�9L&�9��9v�9��9x�9��9'�9�8�9M�9�a�9]s�9��9��9��9}��9���9/��9/��9���9��9���9K��9 ��9���98��9D��98t�9Eb�9xL�9x   x   $�9��9�
�9���9��9
�9��9�$�9�3�9�F�93`�9;z�9��9խ�9���9���9��9��9���9���9r��99��9��9���9ҭ�9��9�y�9�^�9G�94�9x   x   B�9���9��90��9G��96��9�
�9*�9a0�9TK�9�b�9
z�9��9]��9N��9 ��9"��9���9'��9 ��90��9���9���9ӭ�9��9%z�9�c�9
L�90�9��9x   x   D��9y��9}��93��9���9^��9�9��9�0�9pH�9q_�9�y�9���9��9���9���9���9���9e��9���9���9���99��9��9#z�9^�9�G�9�/�9��9u�9x   x   ���9l��9Y��9���9��9?��9��9;�9E)�9}G�95c�9�y�9��9��9��9���9q��9���9���9f��9ؼ�9��9D��9�y�9�c�9�G�9�)�9��94��9���9x   x   a��9���9O��9���9��9��9*�9��9�0�9�K�9x_�9�t�9̓�9n��9���9Q��9?��9;��9���9���92��9]��9=t�9�^�9L�9�/�9��9 �9���9���9x   x   ���9
��9���9���9���9���9=��9��9�/�9G�91a�9$}�9���9U��9��9N��9ױ�9W��9y��9���9���9�|�9>b�9G�90�9��93��9���9��9���9x   x   ���9־�9��9 ��9���9"��9��9,�9/4�9�L�9f�9+y�9��9]��9��9J��9K��9j��9���9���9sy�9�e�9vL�94�9��9p�9���9���9���9���9x   x   ���9���9���9��9��9�)�9A�9�b�9V�9&��98��9���9���9���9]��9���9��9���9Z��9e��9c��9C��9��9Hc�9�@�9@*�9&�9��9���9n��9x   x   ���9���9��9H�9#�9M5�9QU�9Km�9߅�9��9��9���9T��9���9���9
��9���9E��9���9 ��9���9u��9tl�9�V�9�4�9�"�9^�9���9���9���9x   x   ���9���9��9*�9�+�9�E�9;^�9�u�94��9أ�9d��9��9��9S��9{��9���9���9���9���96��9��9�v�9F]�9�D�9�,�9��9��9.��9K��9|��9x   x   ��9B�9"�9`+�90A�9S�9Ti�9z��9+��9��9���9���9���9��9h��9���9���9���9"��9͕�9ҁ�9�i�9�S�9�A�9j)�9j�9��9��9.��9���9x   x   ��9#�9�+�95A�9�W�9�f�9*y�9<��9���9ر�9���9���9t��9��9���9>��9-��9��9:��9i��9�y�9@f�9�V�9�A�9'-�9�!�9v�9<�9�94�9x   x   �)�9D5�9�E�9S�9�f�9�}�9���9��9���9ʹ�9P��9l��9���9���9���9j��9���9���94��9%��9�|�90g�9S�9�D�95�9�+�98)�9x�9� �9�(�9x   x   A�9MU�98^�9Pi�9'y�9���92��9��9s��9ٿ�9��9���9i��9���9���9���9Q��9L��9`��9��9�y�9�h�9�^�9�T�9;A�95A�9^>�9j8�9<=�9eB�9x   x   �b�9Jm�9�u�9u��9<��9��9��9;��9l��9ý�9��9���9���9S��9Ѽ�9ʵ�9���9.��9p��9-��9��98u�9�m�9�c�9�X�9�U�9�U�9�U�9�U�9&Y�9x   x   N�9ׅ�9/��9%��9���9���9q��9b��9���9���9"��9���9r��9���9��9Z��9���9���9���9B��9���9��9R~�9Cx�9�x�9'v�9,s�9Iw�9�v�9`x�9x   x   !��9��9̣�9���9ӱ�9ʹ�9ؿ�9���9���9���9L��9���9=��9
��9���9s��9ȵ�9Q��9��9P��9��9���9��9^��9���9o��9ҏ�9��9���9ɘ�9x   x   3��9׵�9]��9���9���9S��9	��9��9��9F��9g��9R��9���9���9\��90��9ú�9t��9~��9���9Q��9˯�9���9u��93��9��9���9��9s��9���9x   x   ���9���9��9���9���9m��9���9���9���9���9R��9��9���90��9���9���9w��9��9���9���9���9���9���9/��9}��9���9���9!��9o��9���9x   x   ���9H��9��9���9o��9���9k��9���9m��9=��9��9���9(��9y��9���9���9���9��9���9e��9>��9��9���9��9���9Y��9v��9|��9��9-��9x   x   ���9���9M��9��9��9���9���9X��9���9��9���9/��9z��9���9���9���9?��9���9���9���9g�9c	�95�9�9��9 �9	�9W�9� �9	��9x   x   S��9���9u��9d��9���9���9���9Ӽ�9��9 ��9Z��9���9���9���9���9���9���9��9p�9?�9+�9�)�9�)�9�&�9*�9l(�9Y�9��9x�9T�9x   x   ���9
��9���9���9>��9q��9���9ǵ�9b��9x��90��9���9���9���9���9���9q�9��9�#�9�-�9�7�9^C�9E�9�D�9DD�9�7�9&-�9�#�99�9X�9x   x   v��9���9���9���9.��9���9T��9���9���9е�9Ⱥ�9���9��9B��9���9q�9�"�9n0�9�7�9�K�9AQ�9�U�9,^�9sT�95Q�9"K�9�8�9�/�9�"�9|�9x   x   ���9?��9���9���9��9���9P��90��9���9S��9x��9$��9��9���9��9��9t0�98�9~J�97]�9[^�9�f�9Hh�9�^�9y]�9cJ�9�7�9�0�9��9��9x   x   U��9���9���9!��9>��9?��9f��9z��9 ��9&��9���9���9���9���9u�9�#�9�7�9zJ�9S[�9=h�9�r�9_r�9�q�9!h�9l[�9J�9U8�9�#�9/�9���9x   x   e��9���9;��9ʕ�9p��9)��9��95��9E��9b��9���9���9l��9���9@�9�-�9�K�98]�9Dh�9~v�9�x�9�x�9�w�9�g�9�]�9�K�9�,�9��9���9���9x   x   g��9���9��9ׁ�9�y�9�|�9�y�9��9���9��9Y��9���9G��9p�90�9�7�9IQ�9^^�9�r�9�x�9�x�9�x�9r�9g^�9�P�9�7�96�9�9]��9=��9x   x   J��9y��9�v�9�i�9Ef�95g�9�h�9Fu�9��9���9ϯ�9���9��9o	�9�)�9`C�9�U�9�f�9_r�9�x�9�x�9br�9�g�9�U�9�C�9%*�9��9���9^��9T��9x   x   ��9wl�9K]�9�S�9�V�9S�9�^�9�m�9_~�9 ��9���9���9���9?�9*�9E�93^�9Nh�9�q�9�w�9r�9�g�9�\�9~E�9�(�9��9���9���9��9���9x   x   Nc�9�V�9�D�9�A�9�A�9�D�9�T�9�c�9Nx�9g��9���99��9&��9$�9	'�9�D�9�T�9�^�9-h�9�g�9h^�9�U�9}E�9�'�9�9 ��9���9
��9Η�9�x�9x   x   �@�9�4�9�,�9r)�90-�95�9GA�9�X�9�x�9���9A��9���9���9��9*�9KD�9>Q�9z]�9q[�9�]�9�P�9�C�9�(�9�9���9���9��9���9�w�9�W�9x   x   ?*�9�"�9��9v�9�!�9�+�96A�9�U�9,v�9z��9#��9���9d��9�9{(�9�7�90K�9jJ�9 J�9�K�98�9/*�9��9��9���9���96��9�u�9sW�9C�9x   x   )�9b�9��9��9z�9D)�9h>�9�U�92s�9���9���9���9���9	�9b�9--�9�8�9�7�9]8�9 -�97�9��9���9���9��9:��9�s�9�U�9N;�9�)�9x   x   ��9���96��9��9D�9��9w8�9V�9Tw�9&��9'��9)��9���9\�9��9�#�9�/�9�0�9�#�9��9�9���9���9	��9���9�u�9�U�9F:�9� �9�9x   x   ���9���9K��96��9	�9� �9E=�9�U�9�v�9���9���9x��9��9� �9��9B�9�"�9��94�9���9]��9e��9��9ϗ�9�w�9vW�9L;�9� �9��9"��9x   x   u��9���9z��9���9=�9�(�9kB�92Y�9hx�9Ә�9���9��93��9��9\�9[�9�9��9���9���9;��9Z��9��9�x�9�W�9C�9�)�9�9#��9\��9x   x   ��9��9��9[)�9GE�9�a�9���9���9���9��9�	�9�'�9h@�9�S�9+\�9/[�9\�9}P�9�A�9&�9�
�9���9���9���9H��9�`�9-E�9*�9��9p�9x   x   ��9�9O&�9�9�9yP�9�q�9ƍ�9I��9b��9A��9r�9�(�9�8�9$E�9N�9�M�9�G�9s9�9(�9Q�9[��9A��9���9���9�r�9�O�9o9�9�&�9F�9��9x   x   ��9O&�9�8�9�G�9�`�9�z�9���9���9���9���9��9G$�9�3�9�=�9gG�9;�9�2�9z#�9L�9���9��9��9��9"y�9)a�9�H�9�7�9l%�9��9��9x   x   W)�9�9�9�G�9na�9u�95��9���9���9w��9S��9J�9Q$�9.�9�-�91�9�.�9�%�9��9L��91��9k��9���9���9�u�9�_�9�G�9N;�9�(�9�(�9�'�9x   x   BE�9xP�9�`�9u�9ډ�9���9k��9��9���9��9��9U$�9�'�9#�9�%�9�#�9o�9��9	��96��9���9���9��9�u�9�a�9O�9E�9[<�9�>�9�<�9x   x   sa�9�q�9�z�9,��9���9���9n��98��9���9��9��9Z�9a%�9�$�9��9��9��9���9���9n��9���9���9Ԏ�9�y�9�q�9�a�9�X�9�Q�97R�9�W�9x   x   ���9���9���9���9g��9f��9���97��9���9w
�9��9W�9�9��9;�9e�9��9f��9���9j��9ͽ�9��9ӛ�9<��9���9�x�9�r�9�m�9_s�9�y�9x   x   ���9@��9��9���9��97��97��9>��9�	�9��9I�9��9[�9��9�9J	�9��9���9G��9X��9<��9���9U��9D��9��9���9���9P��9ܔ�99��9x   x   ���9Y��9���9s��9���9���9���9�	�9�9��9��9��94�9o�9��9h	�97 �9��9���9���9���9���9Y��9���9D��9M��9���9���9Ҽ�9���9x   x   ��94��9���9Q��9��9��9y
�9��9��9N�9�9��9g�9�9��9�	�9��9��9f��9���9}��9���9���9%��9���9���9���9���9@��9���9x   x   �	�9l�9��9E�9��9��9��9G�9��9��9�9��9��9z�9��9S�9Z�9,�9P�97�9�	�9�9e�9<�95�9�	�9�9��9��9��9x   x   �'�9�(�9C$�9J$�9L$�9U�9Q�9��9��9��9��9��9��9��9u�9x#�9&�9$�9�'�9�%�9�+�9^*�95-�9�+�9t(�9�)�9�+�9y-�9 *�9�*�9x   x   a@�9�8�9�3�9�-�9�'�9c%�9�9\�95�9n�9��9��9w�90$�9y'�9U-�9�2�9�9�9�A�9�E�9�H�9KO�9�S�9MQ�9�S�9P�9nS�9�O�9jI�9�D�9x   x   �S�9E�9�=�9�-�9#�9�$�9��9��9k�9�9}�9��9,$�9�#�9B/�9_>�9DE�9BR�9�]�9�c�9	m�9�t�9�u�9[}�9�}�9\w�9At�9�k�9�d�9�^�9x   x   \�9N�9aG�9�0�9�%�9��9?�9�9��9��9��9y�9t'�9A/�9�E�93N�9�\�9j�9�t�9��9���9���9��9���9e��9��9C��9���9�s�9:i�9x   x   '[�9�M�9�;�9�.�9�#�9��9e�9L	�9m	�9�	�9]�9#�9Z-�9g>�91N�9gZ�9�p�9��9��9u��9��9\��9߰�9��9ư�9`��9i��9���9��9�p�9x   x   \�9�G�9�2�9�%�9m�9��9��9��9< �9��9a�9&�9�2�9IE�9�\�9�p�9*��9ߚ�9���9���9l��9���9R��9���9
��9|��93��9���9��9�p�9x   x   yP�9z9�9{#�9��9��9���9j��9���9��9��97�9$�9�9�9GR�9
j�9��9��9ܲ�9���9���9H��9[��9���9L��9���9���9���9v��9��9aj�9x   x   �A�9�(�9L�9P��9��9���9���9N��9���9m��9P�9�'�9�A�9�]�9�t�9��9���9���9���9���9���9��9���9���9���9���98��9���99t�9�_�9x   x   &�9R�9���98��9:��9t��9w��9`��9���9���9=�9�%�9�E�9�c�9��9~��9��9���9���9���9<��9D��9h��9���9���9���96��9��9�a�9wE�9x   x   �
�9W��9��9r��9��9���9Խ�9E��9���9���9�	�9�+�9�H�9m�9���9"��9p��9M��9���9>��9���9(��9���9���9f��9��9|��9xn�9�I�9b+�9x   x   ���9=��9��9ð�9���9��9��9���9���9���9�9l*�9YO�9�t�9���9c��9���9c��9��9K��9/��9`��9K��9��9��9��9�r�9nN�9R*�9�
�9x   x    ��9���9��9���9��9��9��9h��9h��9���9u�9F-�9�S�9�u�9$��9��9Z��9���9���9l��9���9J��9u��9B��9��9�w�9�U�9�,�9��9���9x   x   ���9���9'y�9�u�9�u�9�y�9H��9R��9���90��9L�9�+�9]Q�9f}�9���9��9���9S��9���9���9���9���9C��9К�9�}�9)N�9�+�9}�9���9��9x   x   M��9�r�93a�9�_�9�a�9r�9���9���9V��9���9F�9|(�9�S�9�}�9s��9а�9��9���9���9���9k��9��9��9�}�9^U�9�)�9Y�9��9;��9���9x   x   �`�9�O�9�H�9�G�9O�9�a�9�x�9ĕ�9]��9���9
�9�)�9P�9iw�9���9i��9���9���9���9���9��9��9�w�9*N�9�)�9k�9,��9i��9���9mz�9x   x   2E�9u9�9�7�9T;�9E�9�X�9�r�9��9��9���9#�9�+�9~S�9Lt�9P��9w��9<��9���9>��9<��9{��9�r�9�U�9�+�9W�9'��9���9���9�p�9�Y�9x   x   
*�9'�9w%�9�(�9e<�9�Q�9�m�9a��9���9���9��9�-�9�O�9�k�9���9���9ę�9}��9���9!��9yn�9nN�9�,�9~�9��9g��9���9�o�9R�9�;�9x   x    �9I�9��9�(�9�>�9?R�9gs�9��9ڼ�9K��9��9*�9}I�9�d�9�s�9���9%��9��9=t�9�a�9�I�9Q*�9��9���95��9���9�p�9R�9X?�9Y(�9x   x   x�9��9��9(�9�<�9�W�9�y�9J��9���9���9��9+�9�D�9�^�9Fi�9�p�9�p�9ej�9�_�9yE�9^+�9�
�9���9��9���9ez�9�Y�9�;�9^(�9��9x   x   �1�9�*�9>�96T�9�o�9���9O��9���9I�9�2�9�`�9��98��9`��95��9���9���9���9��9l��9*a�9�3�9��9g��9���9��9Tp�91U�9r=�9�*�9x   x   �*�9�1�9�H�9�[�9*{�9	��9���9���9��9�;�9@`�9Ѐ�9��9ϯ�9���9���97��9 ��9��9{a�9q:�9��9Z��9x��9%��9�z�94[�9I�9y2�9M)�9x   x   >�9�H�9�[�9Kr�9���9p��9���9���9t#�9�G�9c�9�{�9֏�9ҝ�9���9���90��9|�9�c�9�F�9h#�9���9@��9ŵ�9��9:s�9l[�9�G�9�?�9�6�9x   x   ,T�9�[�9Gr�9���9���9���9���9��9�1�9�I�9Al�9�w�9���9h��9��9r��9Kx�9�k�9lH�9�3�9�9���9}��9f��9���9�q�9�\�98S�9J�9J�9x   x   �o�9!{�9���9���9f��9���9��9�%�9�6�9IS�9�n�9pu�98��9a��9W��9�t�9rn�9�T�9�5�9&�9+�9��9���9��9��9pz�9�p�9�d�9�\�9Fe�9x   x   ���9���9r��9���9���9��9i�9�2�9�G�9�a�9	o�9ou�9z}�9}�9�v�9p�9w`�9�H�9�2�9��9}�9y��9���9w��9��9���9z��9܅�9���9���9x   x   G��9���9���9���9��9m�9O+�9�A�9�V�9�d�9�o�9�s�9�x�9�t�9Xm�9.f�9`V�9�A�9-�9��9��9���9���94��9��9��9��9T��9���93��9x   x   ���9���9���9��9�%�9�2�9�A�9+V�9�a�9�h�9�p�9�y�9@x�9$q�9i�9ab�9?V�9�?�9�2�9&�9z�9,��9��9���9���93��9e��9���92��9H��9x   x   :�9��9p#�9�1�9�6�9�G�9�V�9�a�9�k�9�o�9�m�9Sq�9�m�9-q�9�i�9�a�9�X�9�H�946�9J1�9H%�9	�9��9	�9��9���90��9���93��9x�9x   x   �2�9�;�9�G�9�I�9FS�9�a�9�d�9�h�9�o�9�s�9is�9u�9�q�9�o�9�j�9Jc�9�`�9zS�9XK�9pE�9�:�9�2�9�0�9�/�9f0�9U'�9�'�990�90.�9�1�9x   x   �`�94`�9c�95l�9�n�9o�9�o�9�p�9�m�9hs�93v�9�s�9�o�9�o�9jo�9Lp�9�o�9*j�9�c�9b�9ba�9j`�9�Y�9^\�9P^�9�S�9c]�98]�9�Y�9�`�9x   x   ߁�9ŀ�9�{�9�w�9lu�9nu�9�s�9�y�9Oq�9�t�9�s�9�p�94x�9�s�9v�9�s�9�y�9�|�9�9]�9M��9$��9���9ى�9��9��9��9փ�9��9؃�9x   x   *��9���9ɏ�9y��9,��9u}�9�x�9>x�9�m�9�q�9�o�94x�9�z�94|�9׆�9؅�9���9���9���9*��9��9���9���9���9ϸ�9 ��9Ҳ�9l��9���9��9x   x   U��9Ư�9ʝ�9l��9V��9}�9�t�9%q�9,q�9�o�9�o�9�s�9=|�9H��9w��9���9���9���9��9���9���9���9���9���9���9k��9��9:��9��9���9x   x   2��9���9���9��9S��9�v�9Ym�9i�9�i�9�j�9po�9v�9߆�9p��9��9��9/��9H��9���9y��9���9��9-�9��9t�9�9���9���9���9x��9x   x   ���9���9x��9u��9�t�9p�90f�9cb�9�a�9Sc�9Rp�9�s�9��9���9��9���9���9���9�9��9X&�9�+�95�9|5�9J-�9t&�9��9�9q��9���9x   x   ���94��9+��9Mx�9un�9z`�9hV�9AV�9�X�9�`�9�o�9�y�9���9���95��9���9���9H
�9�"�9K1�9~B�9�O�9�P�9�N�9FB�91�9E"�9	�9%��9=��9x   x   ���9��9�{�9�k�9 U�9�H�9B�9�?�9�H�9�S�9:j�9�|�9���9���9P��9���9J
�9�0�9�D�9�L�9�c�9�g�9�h�9�c�9 M�9�E�9J1�9�9���9���9x   x   ��9��9�c�9jH�9�5�9�2�9-�9�2�9:6�9aK�9�c�9�9���9��9���9�9�"�9�D�9�X�9�k�9
w�9�w�9Qv�9=l�9zW�9cC�9x"�9�9���9���9x   x   f��9a�9�F�9�3�9&�9��9��9%&�9Z1�9{E�9�b�9b�95��9���9���9��9O1�9�L�9�k�9�z�9E��9b��9�z�9�k�9�N�942�9Z�9���9���9���9x   x   (a�9z:�9r#�9�98�9��9��9��9V%�9�:�9sa�9U��9��9���9���9^&�9�B�9�c�9	w�9F��9m��9:��9wv�9Ic�9@�9�'�9��9p��9���9E��9x   x   �3�9��9���9���9��9���9���98��9�9�2�9}`�98��9Ӱ�9���9��9�+�9�O�9�g�9�w�9d��9>��9!x�9�h�9�Q�9M,�9��9���9���9P��9�_�9x   x   ��9^��9E��9���9���9���9���9+��9��9�0�9�Y�9���9��9���9>�95�9�P�9�h�9Vv�9�z�9zv�9�h�9�N�9�5�9��9��9˴�9��9e[�9�0�9x   x   i��9~��9ѵ�9s��9+��9���9F��9��9�9�/�9m\�9��9ĺ�9���9��9�5�9�N�9�c�9Al�9�k�9Pc�9�Q�9�5�9n�9��9q��9���9\�9�.�9|�9x   x   ���9+��9 ��9���9(��9��9��9���9��9u0�9`^�9%��9��9���9��9Y-�9XB�90M�9�W�9�N�9@�9N,�9��9��9��9��90^�9<0�9(��90��9x   x   (��9�z�9Ds�9�q�9�z�9���9+��9C��9���9h'�9�S�9���9.��9~��9*�9&�9	1�9�E�9eC�942�9�'�9��9~��9m��9��9jR�9�(�9P��9)��9h��9x   x   Yp�96[�9u[�9�\�9�p�9}��9��9o��9I��9(�9t]�9+��9��9#��9���9��9Q"�9]1�9�"�9c�9 ��9���9Ѵ�9���92^�9�(�9e��9���9p��9H��9x   x   2U�9I�9�G�9BS�9�d�9��9b��9���9���9I0�9G]�9��9}��9J��9���9'�9%	�9�9�9���9u��9���9��9\�9;0�9M��9���9g��9��9�c�9x   x   y=�9�2�9�?�9J�9]�9ʄ�9���9B��9G��9F.�9�Y�9���9���9��9���9{��9+��9 ��9���9���9���9J��9d[�9�.�9+��9)��9u��9��9�^�9�I�9x   x   �*�9J)�9�6�9 J�9Me�9���9?��9V��9��9�1�9�`�9��9��9���9���9���9I��9���9���9���9I��9�_�9�0�9{�9.��9d��9J��9�c�9�I�9�7�9x   x   <�9�A�9�S�9�h�9��9C��9��9{�9�S�9ǆ�98��9���9U�9� �9$/�9�6�9�-�9Z �9h�9m��9g��9��9�T�9t �9���9/��9���9�i�9�R�9�A�9x   x   �A�9�M�9C[�9�|�9ߡ�9k��9���9i/�9m_�9ŏ�9,��9���9U��9�
�9o�9$�9��9���9��9q��9���9_�9x-�9���9���9��9�z�9�Z�9�N�9[A�9x   x   {S�9C[�9t�9O��9��9���9�9�?�9�j�9���9#��9���9���9���9c�9��9v��9[��9t��9���9fk�9oA�9I�9���9˷�9��9�u�9�Z�9�R�9�I�9x   x   �h�9�|�9O��9Z��9���9o��9j'�9�T�9`{�9��93��9���9���9>��91��9���9���9N��9B��9}�9�R�9�%�9���9c��9���9C��9|�9�h�9�a�9�`�9x   x   ڏ�9ܡ�9��9���9���9�9"@�9�c�9Z��9*��9��9 ��98��9���9c��9���97��9��9��9�c�9�B�9��9v��9%��9��9��9Ӑ�9z��9E�9߂�9x   x   9��9`��9���9n��9�9�C�9�\�9�|�9U��98��9���9	��9��9���9q��9��9���9|��9h}�9g[�9�A�9%�9��9r��9���9��9���9��9ٟ�9���9x   x   ��9{��9�9a'�9@�9�\�9|�9���97��9��9j��9���9���9n��9���9��95��9ƕ�9_|�9�]�9�@�9N&�9�9���9]��9���9,��9l��9���9���9x   x   p�9a/�9�?�9�T�9�c�9�|�9���9���9���9���9k��9?��9$��9���9]��9���9Z��9���9�|�9\c�9U�9�>�9�.�9�9��9
�9� �9� �9�
�9o�9x   x   �S�9\_�9�j�9\{�9T��9U��93��9���9���9��9 ��9���9,��9X��9u��9.��9s��9A��9���9�z�9�l�9_�9�T�9�G�9�<�9`=�9 =�9�;�9�=�9HH�9x   x   ���9���9x��9��9��92��9޹�9���9��9f��9��9��9=��90��9��9T��9g��9��9��9U��9ڎ�9.��9��9z�9&p�9�r�9�t�9�p�9]x�9Ā�9x   x   +��9��9��9-��9��9���9f��9n��9��9��9��9��9)��9���9{��9s��9}��9���9���9%��9%��9:��9��9��9��9X��92��9��9-��9+��9x   x   ���9���9���9���9���9��9���9@��9���9��9!��9���9y��9u��9���9���9���9j��9w��9X��9���9d��9��9+��9���9L��9���9���9���9���9x   x   E�9J��9���9���91��9 ��9���9'��9.��9=��9.��9|��9"��9���9'��9���9���9a��9D�9��9 �9M�9 �9�#�9$�9$�9��9��9��9�9x   x   q �9�
�9���99��9���9���9j��9���9[��93��9���9t��9���9��9���9� �9�
�9� �91.�9>�9�J�9PM�9^V�9�Y�9�X�9W�9NN�9I�9�>�9�/�9x   x   /�9a�9[�9+��9^��9p��9���9^��9|��9��9|��9���9)��9���96�9@�9�.�9{C�9�T�9Fj�9
w�9S��9n��9 ��9Ј�9��9{w�9�j�9�R�9�B�9x   x   �6�9�9��9���9���9��9��9��98��9[��9{��9���9���9� �9E�9?7�9�M�9/h�9��9���9���9ۭ�9���9���9w��9;��9A��9,��9ji�9�M�9x   x   �-�9��9v��9���97��9���98��9\��9}��9n��9���9���9���9�
�9�.�9�M�9�r�9g��9���9���9
��9���9%��9���9��9���9���9���9*r�9�N�9x   x   O �9���9Z��9Q��9��9���9Е�9���9K��9��9���9q��9g��9� �9�C�98h�9j��95��9m��9p��9f��9}��9���9���9���9��9ϩ�9���9�g�9D�9x   x   e�9��9|��9I��9��9s}�9l|�9�|�9ȍ�9��9���9���9S�98.�9�T�9��9���9k��9���9���9��9s�9N�9���9T��9k��9���9 ��9�S�9�.�9x   x   n��9t��9���9#}�9�c�9q[�9�]�9oc�9�z�9d��98��9g��9��9>�9Nj�9ǔ�9���9p��9���9��9v�9�9
�9���9���9l��9���9�k�9C>�9�9x   x   j��9���9hk�9�R�9C�9�A�9�@�9U�9�l�9��97��9���9�9�J�9w�9��9��9m��9��9|�9e�9|�9W�9���9~��9���9�v�9�I�9S�9Z��9x   x   ���9_�9xA�9&�9��95�9c&�9�>�95_�9<��9N��9w��9a�9dM�9]��9��9���9���9t�9�9z�9[�9f��9l��9-��9ǁ�9N�9(�9���9­�9x   x   �T�9~-�9S�9���9���9(��9 �9�.�9�T�9��9��9��91 �9pV�9��9���93��9���9Y�9�9Y�9i��9���98��9ވ�9�V�95�9���9��9��9x   x   � �9���9���9s��94��9���9���9'�9�G�9z�9.��9C��9�#�9�Y�94��9²�9���9���9���9���9���9o��97��9���9EY�9�#�9g��9 ��9y�9(G�9x   x   ���9���9Է�9��9��9���9s��9�9�<�9;p�9���9���9/$�9�X�9ވ�9���9+��9���9`��9���9��93��9߈�9EY�9�$�9���9��9�p�9_>�9��9x   x   2��9!��9��9N��9 ��9)��9���9'
�9t=�9�r�9r��9c��9/$�90W�9��9P��9���9"��9v��9y��9���9Ё�9�V�9�#�9���9���9�s�9�;�9?
�9���9x   x   ���9�z�9�u�9$|�9��9ū�9J��9� �97=�9�t�9I��9���9��9cN�9�w�9U��9���9٩�9���9���9�v�9N�94�9a��9��9�s�9"=�9r�9s��93��9x   x   �i�9�Z�9�Z�9i�9���9��9���9�9�;�9�p�9��9��9��9-I�9�j�9?��9���9��9(��9�k�9�I�9(�9���9��9�p�9�;�9n�9���9Ӡ�9���9x   x   �R�9O�9 S�9�a�9V�9ޟ�9���9�
�9�=�9sx�9D��9���9��9�>�9S�9}i�92r�9�g�9�S�9J>�9X�9���9��9y�9\>�9=
�9k��9Π�9D��9ga�9x   x   �A�9bA�9�I�9�`�9��9���9���9|�9YH�9Ӏ�9?��9���9-�9�/�9�B�9�M�9�N�9$D�9�.�9�9]��9���9���9G�9��9���9,��9���9fa�9J�9x   x   l6�9�C�9�W�9Xu�9r��9O��9	�9�N�9���9?��9�	�9�>�9Dh�9}��9���97��9��9ǒ�9�h�9�=�94	�9���9n��9�O�9A�9m��9Ԡ�9�v�9�U�9{C�9x   x   �C�9�N�9�k�9���99��9��9(-�9�]�9#��9���9j�9=�9e�9�x�9��9��9�w�9�c�9=�9��9q��9��9�]�9�,�9|��9Ƹ�9@��9fk�9�P�9FD�9x   x   �W�9�k�99��9Q��9���9��91B�9�z�9���9���9P�9s8�9ZX�9�f�9Ls�9"h�9�X�9�9�9��9���9���9_{�9LB�9��9���9���9ȇ�96k�9U�9�Q�9x   x   Wu�9��9I��9��9' �9h+�9�g�9]��9%��9���9��9"9�9�L�9/W�9�T�9<L�9�8�9��9���9u��9���9'g�9�+�9[ �9���9U��99��9�v�9�n�9�l�9x   x   h��9-��9���9" �9�)�9	S�9)��9���9���9���92�9r6�9C@�9�I�9nB�9�6�9��9���9��9��9?��9cS�90)�9a �9���9���9��9���9���9V��9x   x   @��9��9~�9a+�9	S�9w�9��9���9z��9��9��9V/�9�?�9�?�9/-�9��9�9���9��9��9�u�9�S�9w+�9��9>��9x��9���9���9ֿ�9���9x   x   ��9-�9$B�9�g�9$��9��9���9��9a��9�9�9�0�9r5�9B1�9U!�9��9P��9���9!��9S��9i��9g�98C�9i,�9��9��99��9n��9T��9Y�9x   x   sN�9�]�9�z�9X��9���9���9��9��9��9� �9D*�9*�9�)�9m)�9��9��9���9���9v��9C��9���9�y�9 ^�9�O�9�A�94�9:3�9w4�9�5�9nA�9x   x   ���9��9���9��9���9t��9^��9��9��9�!�9�*�9�)�9�+�9_!�9'�9B�9j��9a��9��9���9��9͟�9ǌ�9$��9��9v�9�r�9�s�9s�9���9x   x   +��9���9���9���9���9��9�9� �9�!�9f&�9,�9S+�9�&�9�!�9x�9 �9�
�9���9���9���9f��9+��9���9��9���9?��9���9ۿ�9P��9���9x   x   �	�9Z�9A�9��9)�9��9�9@*�9�*�9�,�9�0�9},�9�*�9*�9!�9a�9� �9O�9\�9\�9��9��9��9%�99	�9~
�9�9��9�9�9x   x   �>�9=�9^8�99�9h6�9G/�9�0�9*�9�)�9U+�9},�9!)�9X*�9e2�9�,�9p4�9:�9O9�9�<�9?�9�H�9�F�9�I�9J�9+J�9�J�9�J�9�H�9QG�9	I�9x   x   3h�9�d�9PX�9�L�9B@�9�?�9l5�9�)�9�+�9�&�9�*�9X*�9U3�9�@�9	D�9L�9�W�9;d�9}g�9%w�9�~�91��9_��9B��9^��9y��9���9ͅ�9C~�9�u�9x   x   f��9�x�9�f�9W�9�I�9�?�9A1�9o)�9b!�9�!�9*�9l2�9�@�9�F�9�U�9Eg�9�x�9C��9��9
��9#��9���9���9���9���9���9���9غ�98��9R��9x   x   ���9���9Es�9�T�9oB�9/-�9Z!�9��9%�9x�9/�9�,�9
D�9�U�9�t�9���9 �9���9J��91��9O��9�	�9��9(�9��9��9j��9T��9#��9���9x   x   +��9��9h�98L�9�6�9��9��9��9J�9 �9m�9y4�9L�9Ig�9���9"��9���9B��9%�9��9�,�96D�9H�9�G�91D�9-�9��9 �9���9?��9x   x   Р�9�w�9~X�9�8�9��9�9V��9���9w��9�
�9� �9":�9�W�9�x�9Š�9���9���9��9�7�9O�9a�91t�9|x�9�s�9a�9iO�9�7�9��91��9���9x   x   Œ�9�c�9�9�9��9���9���9���9���9l��9���9X�9c9�9Pd�9T��9���9I��9��9>�9�^�9Vz�9J��9��9���9ȍ�9Ty�9�^�9�=�9��9���9��9x   x   �h�9=�9��9���9#��9#��9-��9���9#��9���9j�9�<�9�g�9��9X��9-�9�7�9�^�9Ƃ�9���9���9���9Z��9C��9.��9d^�9T8�9��9y��9��9x   x   �=�9��9���9}��9 ��9��9c��9U��9���9��9o�9?�91w�9 ��9;��9��9O�9[z�9���9}��9��9���9���9��9�z�9O�9N�9���9��9�v�9x   x   :	�9u��9���9���9N��9�u�9|��9���9��9w��9��9�H�9�~�95��9]��9�,�9a�9P��9���9��90��9)��9��9ی�9�`�9�-�9���9ȹ�9?}�9�I�9x   x   ���9"��9q{�96g�9uS�9�S�9%g�9�y�9��9E��9��9G�9B��9���9�	�9FD�9Dt�9��9���9��9(��9#��9���90u�9C�9��9{��9��9G�9��9x   x   t��9�]�9XB�9�+�9E)�9�+�9RC�9/^�9��9���9�9�I�9{��9���9��9H�9�x�9��9e��9���9���9���9?w�90H�9��9D��9L��9yI�9��9���9x   x   �O�9�,�9��9g �9q �9��9,�9�O�98��9$��9=�9(J�9]��9��9=�9�G�9�s�9֍�9I��9��9��94u�9+H�9�9^��9ԏ�9K�9��9���9��9x   x   I�9���9���9���9���9S��9��9�A�9��9پ�9U	�9CJ�9~��9
��9��9HD�9%a�9dy�97��9�z�9�`�9"C�9��9^��9
��9�I�9��9���9��9=A�9x   x   w��9ϸ�9���9c��9и�9���9��9#4�95v�9_��9�
�9�J�9���9���9 	�9-�9}O�9_�9o^�9O�9�-�9��9D��9؏�9�I�9��9J��9 t�9r4�9��9x   x   ڠ�9H��9҇�9G��9���9���9L��9L3�9�r�9���99�9�J�9ˎ�9���9|��9��98�9�=�9X8�9Y�9���9��9N��9K�9��9F��9Is�9�4�9I��9���9x   x   �v�9ok�9Ek�9�v�9���9���9���9�4�9�s�9���9��9�H�9��9��9j��91�9��9��9��9��9й�9��9vI�9��9���9�s�9�4�9���9O��95��9x   x   �U�9�P�9!U�9�n�9���9��9d��9�5�9��9h��9&�9bG�9Y~�9T��9:��9��9A��9���9���9���9?}�9G�9��9���9��9o4�9I��9M��9u��9Hn�9x   x   �C�9PD�9R�9�l�9h��9���9i�9�A�9���9��9,�9I�9v�9b��9���9H��9���9��9��9�v�9�I�9|�9���9��9?A�9��9���97��9Kn�9cR�9x   x   �1�99�9�O�9/z�9o��9���9/�9���93��9��9�c�9m��9<��9���9��9�&�9��9��9k��9V��9Vb�9��9��9��9�/�9���9/��9U{�93N�9�8�9x   x   9�9�@�9�d�9r��9��9S�9tL�9���9��9N%�9�k�9x��9��9v��9d��9.��9��9^��9���9�l�9�&�9O��9��9�K�9��9���9 ��9Je�9B�9T9�9x   x   �O�9�d�9���9���9���9q*�9p�9���9o��9�8�9�r�9���9i��9k��9��9��9J��9��9�q�9�7�9n��9��9�o�9�*�95��91��9���9�d�9�N�9GJ�9x   x   "z�9i��9���9���9��9�T�9��9���9�9TB�9Rw�9���9���9��9t��9���9ʔ�9�v�9�C�9��9��9���9QU�9�9���9Ѵ�9���9{�9h�9�f�9x   x   f��9��9���9��9bL�9��9׸�97��9W$�9fQ�9#}�9[��9���9���9���9���9�}�9�P�9S$�9K��9d��9���9-K�9l�9%��9���9��9���9���9;��9x   x   ���9A�9k*�9�T�9��9���9K��9��9n9�9�b�9Z�9��9���9h��98��9_�9dc�9f8�9;�9|��9˱�9���9 U�9�*�9��9k��9���9F��9 ��9,��9x   x   	/�9bL�9�o�9ގ�9Ӹ�9M��9]�9$4�9R�9�m�9w��9]��9��9}��9d��9Al�9�S�9�3�9*�9"��9���94��9co�9+L�94/�9�9��9d�9��9��9x   x   ���9���9���9}��91��9��9$4�9�O�9�^�9Dw�9ڄ�9q��9���9 ��9tw�9�^�9�N�95�9y�9���9���9���9M��9c��9Jm�9�_�9,W�9X�9�`�9�m�9x   x   !��9���9b��9�9S$�9c9�9	R�9�^�9_q�9v��9���9n��9���9J��9�r�9w^�92R�9�9�9H#�9%�9���9���9���9?��9���9���9Ŭ�9���9���9Կ�9x   x   ��99%�9�8�9BB�9_Q�9�b�9�m�9?w�9x��99��9!��9|��9���9t��9~v�9�n�9�`�9{R�9�B�9�8�9&�9��9��9�	�9o�9u��9d��9n�9U	�9��9x   x   �c�9�k�9�r�9@w�9}�9R�9z��9ք�9߈�9��9̉�9��9݇�9��9*��9R��9�}�9v�9dr�9_k�9c�9�f�9i_�9._�9[�9�Q�9�X�9_�9J`�9�e�9x   x   T��9g��9���9���9R��9��9d��9m��9n��9x��9��9:��9b��9c��9y��9ݓ�9J��9���9���9��9���9խ�9<��9���9д�9���94��9+��9���9V��9x   x   $��9���9P��9���9��9���9��9���9���9���9߇�9d��9��9���9ݨ�9���9d��9���9���9���9���9���9_�9��9�9��9��9���9���9��9x   x   ���9i��9[��9��9���9a��9���9���9U��9}��9��9`��9���9��9��9<��9���9U��9��90.�9|?�9@L�9GR�9�W�9�W�9�R�9�L�9�=�9e.�9��9x   x   ��9Q��9��9p��9���95��9h��9zw�9�r�9�v�9.��9|��9��9��9���9b��9g�9�8�9�]�9o�94��9ܙ�95��9ͣ�9i��9*��9|��9�p�9'\�99�9x   x   �&�9!��9��9���9���9X�9Gl�9�^�9^�9o�9T��9��9Ʈ�9D��9g��9�'�9JP�9�s�9D��9N��9��9T��9���9U��9k��9���9��9ӕ�9�t�9�O�9x   x   ��9y��9C��9ɔ�9�}�9ic�9�S�9�N�9AR�9a�9�}�9Y��9q��9���9q�9JP�9ʀ�9٤�9���9���90
�9*�9x�9��9�	�9x��9���9���9��9�P�9x   x   ��9T��9��9�v�9�P�9p8�9�3�95�9�9�9�R�9v�9ќ�9���9_��9�8�9�s�9ۤ�9 ��9��9W!�9�>�9�C�9-C�9�>�9� �9��9��9>��9�t�9.8�9x   x   g��9���9�q�9 D�9\$�9H�9@�9��9X#�9�B�9yr�9���9���9��9�]�9R��9 ��9��9/�9�N�9�b�9we�9�b�9cO�9�.�9�9~��9$��9�\�9R�9x   x   Y��9�l�98�9��9^��9���92��9���99�9�8�9zk�9���9���9I.�9)o�9Z��9 ��9a!�9�N�9�i�9ry�9'z�9sh�9SN�9�!�9���9}��9>o�9a1�9
��9x   x   Tb�9�&�9y��9��9w��9߱�9���9���9��9$&�9:c�9��9���9�?�9M��9��9?
�9�>�9�b�9uy�9ׄ�9�y�9�c�9�>�9�
�9��9���9�<�9���9���9x   x   ��9U��9���9���9���9͆�9J��9���9���9�9�f�9���9���9YL�9���9e��9>�9�C�9�e�9*z�9�y�9e�9$C�9/�9��9���9EN�96�9P��9�f�9x   x   "��9��9�o�9fU�9HK�9U�9o�9o��9���9��9�_�9[��9�9aR�9P��9���9��9?C�9�b�9yh�9�c�9 C�9��9<��9p��9�Q�9�9#��9_�9��9x   x    ��9�K�9�*�9&�9��9�*�9ML�9���9Y��9�	�9P_�9���9��9�W�9��9n��9��9�>�9sO�9`N�9�>�93�9;��9��9�W�9}�9d��9f`�9	�9���9x   x   �/�9��9I��9���9<��9��9R/�9pm�9���9��9)[�9���9;�9X�9���9���9�	�9!�9�.�9�!�9�
�9(��9w��9�W�9
�9��9eY�9��9���9�m�9x   x   ���9���9C��9��9���9���9�9�_�9���9���9�Q�9ĵ�9��9�R�9K��9���9���9��9�9���9��9���9�Q�9{�9��9(S�9���9î�9_�9��9x   x   ;��9��9��9���9���9���9��9KW�9��9���9Y�9X��9��9�L�9���9��9���9��9���9���9���9IN�9�9e��9bY�9���9��9oX�9��9H��9x   x   ^{�9Se�9�d�9!{�9���9d��9��95X�9���9��99_�9L��9���9>�9�p�9��9���9M��9-��9Ao�9�<�9;�9"��9f`�9��9Ʈ�9nX�9��9g��9ՙ�9x   x   9N�9B�9�N�9#h�9
��9��9��9�`�9س�9v	�9i`�9̭�9��9z.�9?\�9�t�9��9�t�9�\�9a1�9���9S��9_�9	�9���9_�9��9a��9��9�g�9x   x   �8�9X9�9VJ�9�f�9G��9B��9��9�m�9��9��9f�9o��9#��9��929�9�O�9�P�9;8�9\�9��9���9�f�9��9���9�m�9��9G��9͙�9�g�9pK�9x   x   ��9��9�0�9/^�9ƞ�99��9�J�9 ��9��9�e�9���9!�9�S�9F��9��9���9���9��9�S�9�9���9�e�9 �9��95L�9���9x��9�^�9�0�9��9x   x   ��9l+�9%K�9�~�9���9�9�e�9���9J�9�t�9���9��9�=�9�b�9�v�9#w�93a�9�;�9��9���9�u�9��9w��9)e�9��9��9p}�9
L�9�*�9��9x   x   �0�9+K�9u�9x��9g��9�?�9ő�9��9;�9f��9���9��9�-�9�K�9�R�9_L�9d/�9�9���9ց�9�9�9g��9���9�?�9B��9���9�t�9eK�9�1�9�&�9x   x   ^�9�~�9w��9r��9�*�9�s�9���9��9DX�9��9���9'�9�!�9�-�9;-�9�!�9� �9��9���9YW�9��9!��9�t�9�*�9���9Z��9u}�9$^�9�S�9�S�9x   x   ���9���9]��9�*�9ud�9v��9���9�0�9�r�9.��9���9���9�9��9��9���9���9���9{s�9�/�9���9���9&c�9�+�9?��9���9��9}��9n��9���9x   x   $��9	�9�?�9�s�9l��9���9��9Z�9��9��9H��9���9��9w�9��9���9'��9���9�Z�9��9��9���9�s�9u@�9��9���9���9��9'��9}��9x   x   �J�9�e�9���9v��9���9��9UN�9	��9��9W��9*��9���9���9,��9g��9���9~��9X�9[N�9H�9���9���9ޏ�9sf�9�K�9�/�9��94�9V!�9/�9x   x   ��9ܿ�9���9��9�0�9Z�9
��9���9���9���9%��9���9���9F��9���9��9���9���9�Y�9N2�9��9���9���9P��9��9���9Ew�9+w�9���9T��9x   x   l�9/�9;�92X�9�r�9��9��9���9��9���9*��9���9��9l��9\��9���9��9���9�q�9�X�9	9�9.�9��9y��9T��9���9'��9���9���9{��9x   x   ge�9~t�9R��9��9#��9��9O��9���9���9���9|��9���9��9'��9d��9{��9���9��9���9΂�9�u�9Vd�9�X�9SQ�9"E�9�J�9�K�9EE�9�P�9�X�9x   x   ���9h��9��9���9���9?��9$��9��9.��9x��9���9e��9���9K��9P��9���9(��9
��9<��90��9���9��9Y��9���9p��9���9��9!��9��9Q��9x   x   	�9��9��9�9���9���9���9���9���9���9j��9��9���9���9%��9���9� �9�9��9Q�9"
�9N�9G�9��9'�9��9��9�9�9C
�9x   x   jS�9s=�9�-�9�!�9��9��9��9���9��9��9���9���9A��9K�9��9�"�9T.�9P<�9#T�9b[�9k�9�x�9M�9���9i��9���9�~�92z�9l�9�[�9x   x   )��9�b�9�K�9�-�9��9u�9-��9D��9j��9!��9O��9���9T�9��9%.�9#K�9�b�9���9��9���9���9���9���9���9K��9���9���9^��9���9���9x   x   ���9�v�9~R�93-�9��9��9f��9���9`��9o��9Y��9.��9��9 .�9�Q�9�w�9p��9U��9U��9��9q"�9�4�9�J�9�I�9RI�9�4�9�"�9�99��9��9x   x   ���9w�9TL�9�!�9���9���9���9��9���9���9���9���9�"�9&K�9�w�9=��9?��9�	�9�5�9�[�9�t�9���9Ϙ�9���9��9�u�9Z�9�4�9��9��9x   x   ���90a�9f/�9� �9���9/��9���9Ο�9���9��9=��9� �9f.�9�b�9y��9E��9��9�N�9�z�9m��9O��94��9a��9���9��9���9�{�9MP�9��9x��9x   x   ؄�9�;�9�9��9���9���9g�9���9���9$��9��9�9^<�9���9a��9�	�9�N�9*��9���9J��9��9��9�9�9���9x��9g��9N�9�9��9x   x   �S�9��9���9���9�s�9�Z�9kN�9�Y�9�q�9���9Z��9�9?T�9���9a��9�5�9�z�9���9���9��9�-�9I;�9#/�9]�9���9���9�|�984�9��9%��9x   x   �9���9ځ�9fW�90�9��9Y�9h2�9�X�9��9I��9i�9�[�9��9�9�[�9{��9Q��9��9�<�9�M�9N�9�:�9��9���9N��9�[�9��9p��9�Z�9x   x   ���9�u�9�9�9��9���94��9���9��9*9�9�u�9���9F
�9k�9���9�"�9u�9d��9��9�-�9�M�9}R�9�M�9�/�9T�9E��91u�9�#�9{��95k�9��9x   x   �e�9��9y��9;��9���9��9���9���9S�9{d�9��9y�9�x�9��9�4�9���9F��9��9W;�9$N�9�M�9�:�9F�9.��9Ӆ�9�2�9E��9�z�9�9J��9x   x   #�9���9���9�t�9>c�9�s�9���9���9�9�X�9y��9i�9q�9���9�J�9��9}��9(�93/�9�:�9�/�9B�9���9���9�K�9���9�}�9��9���9Y�9x   x   '��97e�9�?�9�*�9�+�9�@�9�f�9u��9���9�Q�9Ȳ�9��9Ɔ�9���9J�9���9���9*�9o�9��9]�95��9���9"J�9&��9���9I�9#��9=P�9d��9x   x   9L�9��9W��9���9Z��9��9�K�92��9x��9ME�9���9J�9���9w��9pI�9-��90��9���9���9���9K��9ׅ�9�K�9$��9P��9��9,��9�D�9���9X��9x   x   ���9��9��9t��9���9���9�/�9���9���9�J�9���9��9τ�9���9�4�9�u�9��9���9���9`��9:u�9�2�9���9���9��9P��9�K�9>��9Q��9j.�9x   x   ���9�}�9�t�9�}�9��9���9��9nw�9Q��9�K�9@��9��9�~�9���9�"�9"Z�9�{�9{��9}�9�[�9�#�9G��9�}�9J�90��9�K�9 ��9	x�91#�90��9x   x   �^�9L�9oK�99^�9���91��9O�9Mw�9��9nE�9G��97�9Vz�9��9?�9�4�9dP�9N�9L4�9��9���9�z�9��9��9�D�9=��9�w�9��9���9���9x   x   �0�9�*�9�1�9�S�9���9>��9r!�9х�9���9�P�9?��9H�93l�9���9Z��9	�9��9�9*��9��9@k�9�9���99P�9���9N��9*#�9���9���9S�9x   x   ��9��9�&�9�S�9���9���9=/�9p��9���9�X�9p��9d
�9�[�9���9��9��9���9"��9*��9�Z�9��9>��9Y�9a��9M��9b.�9-��9���9S�9�'�9x   x   	��9g��9��9�5�9���9��9PO�9���9�:�9V��9��9�w�9)��9��9�.�9&9�9�/�9V	�9L��9Ny�9h�9��9�8�9���9 P�9���9G��9�5�9��9���9x   x   ]��9��9A�9�^�9���9��9�z�9���9CV�9N��9�"�9`v�9Ӹ�9u��9���9���9���9��92v�9�!�9���9�V�9���9${�9t�9:��9�^�9T�9���9q��9x   x    ��9B�9�M�9D��9���9D�9@��9��9�r�9���9�*�9{p�9��9	��9���9'��9_��9�p�9U*�9���9�q�9�9��9�C�9'��9{��9tM�9�9���97��9x   x   w5�9�^�9:��9G��9�+�9�~�9O��9�<�97��99��9�+�9�h�9=��9��9��9e��9�f�9�,�9���9���9�?�9���9��9E+�9���9���9�]�9=6�9#�9�#�9x   x   ���9���9���9�+�9�v�9���9F�9�i�9��9� �9�9�9e�9:z�9s��9�y�9qe�9/:�9) �9Y��9ui�9�9`��9v�9�,�9���9��99��9ch�9�\�9�h�9x   x   i��9��9D�9�~�9���9�9�Z�9���9���96�9�B�9�V�9�o�9so�9�V�9�B�9\�9���9%��9�[�9a�9���9�~�9�D�9p�9N��9i��9y��9Z��9���9x   x   3O�9�z�9&��9B��9;�9�Z�9���9��9���9d'�9�C�9�U�9�]�9�V�9"C�9 &�9���9���9��9�Y�9��9���9>��9c|�9]O�9<,�9v�9��9��9J,�9x   x   ���9���9��9�<�9�i�9���9��9���9��95�9�R�9XT�9�S�9R�9L7�9��9(��9���9���9k�9�<�9��9���9���9R��9���9$��9���9��9'��9x   x   :�9&V�9�r�9 ��9յ�9���9���9��9�-�9RC�9�S�9�R�9�T�9bB�9,�9��9��9���9ҵ�9r��9�p�9�V�92:�9l#�9�9��9 ��98�9*�9�"�9x   x   1��93��9���9#��9� �90�9Z'�95�9NC�9NK�9HR�9�P�9L�9�C�9�5�9P'�9��93�9���9���9q��9���9���9m��9���9��9���9��9]��9���9x   x   ��9~"�9�*�9�+�9�9�9�B�9�C�9�R�9�S�9FR�9 W�9=R�9�R�9S�9�B�9�A�9�8�9.-�9�*�9!�9��9��9T�9��9��9��9^�9H�9��9��9x   x   cw�97v�9]p�9ph�9e�9�V�9�U�9\T�9�R�9�P�9;R�93S�9�T�9�U�9pX�9�f�9�f�9zp�9+v�9vx�9���9���9���9���9���9m��9���9M��9��9��9x   x   ��9���9ӟ�9(��93z�9�o�9�]�9�S�9�T�9L�9�R�9�T�9�]�9�o�9Vv�9���9���9���96��9���9���9���93
�9U�9a�9�	�93
�9���9���9��9x   x   ��9[��9���9ȟ�9k��9po�9�V�9R�9lB�9�C�9!S�9�U�9�o�9��9���9���9���9��9�"�9�E�9Y^�9�t�9��9x��9��9P��9At�9�]�9�D�9�"�9x   x   w.�9���9���9��9�y�9�V�9$C�9U7�9�,�96�9�B�9vX�9]v�9͠�9���9���9V/�9�^�9��9��9 ��9���9���9��9���9H��9���9α�9���9i_�9x   x   9�9���9��9_��9pe�9 C�9"&�9��9��9X'�9�A�9�f�9���9���9���97�9ux�9O��9���9��9E2�9oS�9?Y�9Y�9�S�9�2�9;�9q��9���9�x�9x   x   �/�9���9X��9�f�93:�9f�9���9;��9"��9��9�8�9�f�9���9���9]/�9wx�9���9���9b<�9�i�9��9���92��9��9���9j�9�=�9��9���9�v�9x   x   J	�9
��9�p�9�,�92 �9���9���9���9���9J�9H-�9�p�9���9��9_�9W��9���9AJ�9��9e��9���9���9���9���9۹�9d��9�H�9
��9���9�]�9x   x   H��9/v�9U*�9���9e��9<��9%��9���9��9��9�*�9Pv�9N��9 #�9���9���9p<�9��9���9���9v�9k�9��9W��9v��9J��9V>�9���9`��95#�9x   x   Fy�9�!�9���9���9�i�9�[�9�Y�96k�9���9��9;!�9�x�9���9"F�9
��9��9�i�9p��9���9-)�9�8�9h9�9�'�9���9l��9�g�9��9J��9KF�9��9x   x   h�9���9�q�9�?�9�9��9��9�<�9)q�9���9��9ۈ�9���9�^�9��9]2�9��9���9��9�8�9{C�9%9�9L�9���9���9V1�9���9�]�9B��9j��9x   x   #��9�V�9�9��9��9���9���9��9	W�9���9��9ߊ�9���9 u�9	��9�S�9̨�9���9w�9p9�9'9�9��9O��9��9U�9���9u�9���9��9:�9x   x   �8�9���9��9��9)v�9�~�9f��9��9b:�9���9��9���9`
�9��9��9_Y�9P��9��9��9�'�9W�9R��9%��9"X�9w��92��9[
�9��9��9��9x   x   ���9<{�9�C�9b+�9�,�9�D�9�|�9��9�#�9���9��9ʐ�9��9���95��9CY�9%��9���9k��9���9���9���9'X�9n��9��9m�9̐�9��9J��9*%�9x   x   P�9��9B��9��9���9��9�O�9���9;�9ō�9��9Î�9��9G��9���9�S�9֒�9���9���9x��9���9U�9{��9��9=�9���9i�9���9k�9Ǥ�9x   x   ���9F��9���9���9
��9u��9f,�9	��9,�9V��9$	�9���9'
�9���9t��93�95j�9���9c��9�g�9h1�9���97��9l�9��9:	�9Ҁ�9��9ܐ�9�+�9x   x   W��9�^�9�M�9�]�9Z��9���9��9O��9M��9ƀ�9��9*��9f
�9ot�9���9V�9�=�9�H�9e>�9��9���9u�9^
�9ʐ�9h�9̀�9���9O��9,�9���9x   x   �5�9e�9+�9Y6�9�h�9���9��9Ê�9j�9��9z�9���9��9^�9���9���96��9,��9���9V��9�]�9���9��9��9���9��9O��9}�9���9wh�9x   x   ��9���9��98#�9�\�9���9�9��9W�9���9��9��9���9�D�9���9ۮ�9���9���9j��9SF�9B��9��9��9I��9c�9ݐ�9.�9���9?^�9�"�9x   x   {��9w��9A��9�#�9�h�9��9k,�9N��9�"�9��9��9/��9>��9�"�9�_�9�x�9�v�9^�9<#�9 ��9p��96�9��9%�9���9�+�9���9rh�9�"�9n��9x   x   �d�9Sx�9ƣ�9��9�K�9i��9xC�9���9	c�9���9n�9v��9�N�9E��9ȿ�9���9��9��9KN�90��9n�9���9 b�9"��9�B�9���9�L�9i��9���9�x�9x   x   Nx�9��9���9�9}~�9���9�t�9���9��9#�9@�9���9�4�92t�9k��9E��9t�9�5�9��9~�9.�9��9��9�u�9���9{}�9��9{��9���9�z�9x   x   ���9���9�9�^�9W��9�4�9M��9i0�9��9 �9V��9���9��9�F�9 O�9(F�9� �9��9���9>"�9R��9�.�9��9�4�9L��9`^�9��9���9ġ�9z��9x   x   ���9�9�^�9V��9�9���9k��9<f�9��9�<�9I��9y��9=�9��9��9�9���9��9�;�9���9�g�9.��9���9��9��90^�9��9���9���9��9x   x   �K�9k~�9O��9��9Pv�9~��9C<�9.��9��9<U�9���9���9���9���9:��9���9��9T�9+�9m��9�9�9���9�v�9��9W��9��9�I�9�,�9L#�9|,�9x   x   D��9���9�4�9���9{��9{+�9��9h��9�'�9sk�9��9/��9���9���9���9��9Sl�9�'�9��9���9O-�9#��9C��9�4�9S��9���9(��9���9G��9��9x   x   PC�9�t�94��9U��95<�9��9"��9�9�S�9���9���9���9��9=��9���9g��9�S�9�95��9Q��9�<�9���9��9pv�9�A�9�%�9��9���9��9&�9x   x   ���9���9J0�9%f�9��9a��9�9<N�9Qu�9h��9��9&��9���9���9@��9�t�9|N�9��9���9Q��9�e�9�0�9���9f��9��9��9���9b��9z��9~��9x   x   �b�9݇�9̫�9���9��9�'�9�S�9Qu�9y��9"��9���91��9y��9���9���9�u�9HR�9�&�9�9���9��9'��9`a�9#D�9�1�9!'�9�(�9�'�9�1�9D�9x   x   ���9��9��9r<�9'U�9ek�9���9b��9��9��9��93��9&��9��9��9(��9�m�9�T�9�:�9�!�9��9%��9���9���9���9��9���9���9m��9���9x   x   �m�9�9;��91��9���9��9���9��9���9��9��9��9���9_��9���9E��9W��9���9��9+~�9�m�9�n�9)j�9�_�9�a�9|\�9kb�9L`�9j�9!o�9x   x   J��9���9���9a��9���9��9���9"��91��9;��9��9��9���9"��9���9^��9B��9���9���97��9���9���9���9�9��9��9��9��9s��9��9x   x   �N�9�4�9��9*�9���9���9��9���9z��9-��9���9���9���9'��9I��9��9Y �96�9jM�9/g�9�v�9��9���9��9@��9ܟ�94��9���9�t�9�h�9x   x   !��9t�9�F�9��9���9���9<��9���9���9��9f��9)��9+��9� �9�9TF�98s�9���9���9���9I�9�"�9D,�9�=�9�=�96+�9�!�9�9���9o��9x   x   ���9J��9O�9��93��9���9���9D��9���9���9���9���9O��9�9uN�9��9#��9o��97�9�`�9i��9���9���9p��9��9��9���9xa�9�7�92��9x   x   ���91��9F�9�9���9��9u��9�t�9�u�9=��9Z��9q��9��9^F�9���9���9��9c�9 ��9P��9�9,�9�=�9�=�9�*�95�9��9���9�c�9o�9x   x   ��9t�9� �9���9��9\l�9T�9�N�9_R�9�m�9j��9b��9i �9Fs�93��9��9�z�9K��9f�9�O�9�{�97��92��9���9�{�9XP�9��9���9ry�9��9x   x   ْ�9�5�9���9��9*T�9�'�9.�9�9�&�9�T�9���9���966�9ғ�9���9c�9R��9u#�9�r�9���9��9���9���9o��9��9�q�9�"�99��9�e�9@��9x   x   >N�9��9��9�;�99�9��9R��9���9/�9�:�99��9���9�M�9���9%7�99��9q�9�r�9��9���9f$�9b-�9�$�9���9���9�s�9��9���9)6�9���9x   x   5��9%~�9J"�9���9���9���9r��9}��9���9"�9Y~�9j��9]g�9���9�`�9n��9�O�9���9���9�,�9pK�9�K�9�,�9X��9��9AO�9��9ra�9���9�f�9x   x   n�98�9_��9�g�9�9�9m-�9�<�9f�9:��9,�9n�9���9�v�9r�9���96�9�{�9��9p$�9yK�9 d�9�K�9"%�9���9~�9S�9���9�9�v�9���9x   x   ���9��9/�9L��9���9H��9��9�0�9X��9Y��9%o�9��9J��9�"�9���9?,�9W��9���9u-�9�K�9�K�9�,�9I��9h��9�,�9���9"�9��9���9^o�9x   x   b�9�98��9ԁ�9w�9s��9K��9!��9�a�9���9nj�9!��9���9u,�9ѹ�9�=�9T��9���9�$�9�,�9-%�9C��9x��9�=�9���9�+�9���9���9�i�9���9x   x   .��9v�9	5�9��9�9�4�9�v�9���9ZD�9���9;`�9B�9L��9�=�9���9>�9��9���9���9o��9���9j��9�=�9#��9�=�9j��9��9p`�9W��9NE�9x   x   �B�9���9l��9��9}��9���9�A�9B��9�1�9)��9�a�9��9z��9�=�9C��9+�9�{�9!��9���9 ��9~�9�,�9���9�=�9#��90�9�b�9���9B0�9Q��9x   x   ���9�}�9^�9S^�9!��9���9&�9F��9^'�9R��9�\�9��9��9i+�9��9f�9}P�9�q�9�s�9YO�9b�9���9,�9m��9.�9�\�9���9�)�9���9z&�9x   x   �L�9��9�9��9J�9a��9&	�9���9)�9=��9�b�9��9p��9,"�9̉�9K��9��9�"�9��9#��9ŉ�9"�9ś�9��9�b�9���9�'�9���9	�9��9x   x   v��9���9���9���9�,�9ҋ�9��9���9�'�9(��9�`�9F��9���9>�9�a�9Ţ�9��9Y��9���9�a�9�9��9���9l`�9���9�)�9���9���9��9�,�9x   x   ���9��9��9��9m#�9o��9��9���9�1�9���9Pj�9���9,u�9���9�7�9�c�9�y�9�e�9>6�9���9�v�9���9�i�9R��9;0�9���9	�9܋�90$�9��9x   x   �x�9�z�9���9'��9�,�9I��9*&�9���9>D�9 ��9Uo�9N��9�h�9���9[��9��9��9Y��9���9�f�9���9co�9���9EE�9G��9i&�9��9|,�9���9	��9x   x   ���9��9/(�9��9:��9[��9�#�9���9��9F0�9^��9�e�9���9;�9�m�9���9o�9�8�9���9�f�9>��941�9��9L��9v"�95��9���9�~�9�*�9A��9x   x   ���9��9DY�9���9�2�9���9y^�9��9ݦ�9�M�9p��9�V�9ȷ�9=�9k&�9>%�9� �9��9PW�9{��9�L�90��9x�9B_�9���9l2�9y��9�W�9j�9H��9x   x   '(�9@Y�9���9��9r��97�9��9!D�9@��9�d�9���9�S�9��9��9���9��9ќ�9�Q�9���9vf�9|��9�C�9ߩ�9��9ą�9��9+��9JZ�9�'�9#�9x   x   ��9��9��9�n�9���9[s�9'��9%��9Z�9Ո�9���9K�9ǃ�95��9$��9��9}K�9���9���9g�99��9���9/s�9���9p�9+�9i��9|��9�`�9Ia�9x   x   ��9�2�9]��9���9[�9T��9hV�9a��9�B�9,��9��9<�9jg�9r�9Kg�9e=�9H �9ڭ�9FE�9$��9�T�9��9Y\�9���9m��9�3�9���9���95��9^��9x   x   :��9���9"�9Gs�9K��9�I�9���9��9\{�9m��96
�9�;�9P�9�P�9�:�95	�9���9J{�9��9���9rJ�9���9t�9!�9���9s��9P�90B�9�C�9~P�9x   x   v#�9T^�9���9��9`V�9���9��9�^�9E��9���9<�9%5�9�A�9�4�9�9���9>��9b_�9d�9g��9�W�9���9���9q_�9"�9���9!��97��92��9���9x   x   ���9��9D�9��9K��9��9�^�9Θ�9���9>�9��9�/�9w/�9��95�9���9��9_�9��9���9��9wD�9� �9���9���9i��9�w�9�w�9@��9~��9x   x   b�9���9��9>�9�B�9P{�9C��9���9v��9��9q$�90�9�$�9M�9- �9���98��9�z�9�D�9��9���9���9�~�9�`�9mF�9�1�9P*�92�9F�9�`�9x   x   0�9�M�9�d�9���9��9^��9���98�9��9C&�9�,�9�,�9A&�9P�9"�9L��9l��9��9���98f�9�L�9�0�9�9e�9N��94��9���9)��9�9�9x   x   &��9:��9���9���9l�9*
�94�9��9r$�9�,�9+�9�,�9�$�9x�9�9��9Q �91��97��9���9}��9i��9G��9��9~��9��9��9���9��9���9x   x   �e�9�V�9�S�9�J�9�;�9�;�95�9�/�90�9�,�9�,�9 0�90/�9�3�9�;�9�=�9�J�9(R�9�V�9�f�9�h�9As�9�z�9�9���9Ѓ�9F}�9�z�9t�9ci�9x   x   ���9���9��9���9Ug�9P�9�A�9y/�9�$�9F&�9�$�9:/�9C�9P�9g�9���9Ӝ�9���9���9���9+�9,�9�2�9
?�9;�9�A�9�2�9�+�9w�9O��9x   x   �:�9�9���9#��9�q�9�P�9�4�9��9W�9U�9��9�3�9$P�9{r�9���9k��9* �9]9�9Qi�9���9��9���9���9���9���9���9%��9N��9Y��9�g�9x   x   ~m�9E&�9���9��9@g�9;�9�9A�9? �94�9�9�;�9g�9���9��9{%�9�n�9Y��9��9�0�97_�9 ��9
��9֢�9`��9.��9L^�9�/�9���9���9x   x   ���9 %�9��9ۂ�9e=�9>	�9���9���9���9c��9��9�=�9���9v��9�%�9��9M��9:1�9���9���9� �9� �9�4�9�5�9R�9���9���9Ԃ�9 2�9���9x   x   �n�9� �9Ȝ�9}K�9K �9��9R��9���9N��9���9i �9�J�9��9; �9�n�9V��9sE�9��9�9�M�9E��9~��9t��9��9|��9�M�9�9���9�C�94��9x   x   �8�9 ��9�Q�9���9��9]{�9�_�97_�9 {�9?��9P��9NR�9ݹ�9{9�9n��9L1�9��9��9�w�92��9��9g�9p�9*��9���9�v�9i�9��942�9��9x   x   ���9MW�9���9���9_E�9��9��9��9�D�9Ї�9o��9�V�9���9}i�9.��9Ӄ�9)�9�w�9^��9�"�9�Q�9,]�9R�9�!�9
��9x�9L�9z��9k��9j�9x   x   �f�9u��9�f�9|�9?��9��9���9���9��9nf�9$��9�f�9���9���9�0�9��9�M�9H��9�"�9�c�9���9҃�9�d�9�"�9d��9O�9���9�0�9���9E��9x   x   F��9�L�9���9S��9U�9�J�9�W�9K��9��9�L�9���9"i�9a�9;��9d_�9� �9h��93��9�Q�9Ą�9ƕ�9���9Q�99��9h��9���9�]�9���9��9�h�9x   x   I1�9I��9�C�9���9B��9��9���9�D�9��9�0�9���9�s�9X,�9���93��9� �9���9��9C]�9���9���9c]�9��9}��9��9"��9��9�+�9�t�9u��9x   x   ��9��9��9Ws�9�\�9Ot�9��9� �9�9^�9���9�z�9�2�9��9A��9�4�9���9��94R�9�d�9Q�9��9���9�5�9ќ�9���9�3�99{�9���9u�9x   x   g��9Z_�9��9���9���9\�9�_�9���9�`�9��9a��9R�9X?�9��9��9�5�9Q��9Q��9�!�9�"�9K��9���9�5�9n��9G��9{@�9�~�9���9�	�9�`�9x   x   �"�9���9��97p�9���9��9O"�9E��9�F�9���9ѻ�9ԅ�9V;�9/��9���9��9���9��9+��9}��9}��9��9Ҝ�9H��9�;�9l��9���9���9]E�9'��9x   x   N��9�2�9
�9Z�94�9���9!��9���9�1�9���9;�9��9/B�92��9p��9���9�M�9�v�9/x�9"O�9���90��9���9~@�9o��9��9���93�9 ��9��9x   x   ���9���9L��9���9���9RP�9]��9Bx�9�*�9!��9f��9�}�9J3�9i��9�^�9���9>�9��9j�9���9^�9!��9�3�9�~�9���9���9+�9lw�9���9RP�9x   x   �~�9X�9mZ�9���9���9jB�9q��9�w�9T2�9p��93��96{�9<,�9���9�/�9��9!��95��9���9�0�9���9�+�9<{�9���9���93�9gw�9���9�B�9���9x   x   �*�9x�9�'�9�`�9d��9�C�9k��9���9^F�9P�9U��9`t�9��9���9��9R2�9�C�9T2�9���9���9��9�t�9���9�	�9UE�9��9���9�B�90��9>a�9x   x   Q��9W��99�9ha�9���9�P�9���9���90a�9M�9���9�i�9���9�g�9���9���9X��9���9"j�9J��9�h�9n��9p�9�`�9��9��9EP�9���99a�9'�9x   x   �(�9�9�9#y�9c��9}�9_$�9���9���9ۚ�9�g�9Q-�9���9]t�9���9�"�9�8�9�$�9���9�r�9���9�.�9Uh�9!��9���9���9�%�9�z�9���9e{�9:�9x   x   �9�9�a�9B��9+�9p��9q�9�3�9P�9��9���9s:�9���90S�9���9u��9D��90��9�U�9���90:�9���9}��9B �9U3�9dp�9���9y-�9��9J`�9O8�9x   x   y�96��9�9<��9x"�95��9ׇ�9�H�9$�9��9�O�9���9t+�9ag�9���9�i�9�*�9&��9%P�9t��92�9 I�9ڈ�9��9�!�9 ��9��9���9|�9�j�9x   x   G��9�*�91��9��9P��9�D�9���9w��9aC�9_��9�Q�9t��9s�9�/�9�.�9J
�9���99S�9���9�B�9U��9���9NC�9n��9!�9=��9D,�9	��9���9���9x   x   �|�9Q��9h"�9N��9%.�9M��9�^�9��9W��9M��9;k�9���9]��9��98��9ƺ�9j�96��9���9���9W_�9���94/�9��9P"�9���9,}�9*K�9�1�9I�9x   x   0$�9�p�9��9�D�9E��9�G�9c��9uQ�9���9�&�9�~�9��9���9���9���9f}�9c(�9j��9tO�9��9�F�9���9<E�9i��9q�9�#�9%��9���9	��9���9x   x   ���9�3�9���9���9�^�9_��9|B�9���9a��9"H�9P��9���9���9���9Y��9vI�9]��9\��9D�9=��9�_�9���9��9{3�9���9d��9M��9Y��9'��9i��9x   x   |��9�9YH�9U��9���9lQ�9���9���9�5�9�l�9!��9h��9٥�9��9�j�9�5�9!��9{��9�P�98��9���9I�9W �9ֻ�9u��9Zi�9HX�9�W�9i�9c��9x   x   ���9���9��9;C�9?��9���9Q��9�5�9/Z�9���9���9���9A��9�9�[�9�6�9O��9��9ڄ�9�B�9��9���9&��9�j�9�L�9;�9�0�9%<�97M�9�j�9x   x   �g�9~��9��9<��9/��9�&�9H�9�l�9���9��9���9g��9	��9݆�9Bj�9�G�9:)�9��9���9���9��9
g�9�I�9�3�9K(�9��9z�9'�9 4�9�J�9x   x   -�9>:�9�O�9zQ�9k�9�~�9A��9��9���9���9¦�9���9���9 ��9n��9�|�9jj�9=S�9O�9L:�9U.�9"�9X�9��9��9��9��9Q�9��9~"�9x   x   ]��9���9T��9P��9v��9ݯ�9��9g��9���9k��9���9U��9��9s��9-��9��9���9���9<��9 ��9���9R��9n��9��9��9�9�9���9k��9,��9x   x   "t�9S�9M+�9O�9A��9���9���9ե�9>��9��9���9��9
��9!��9��9O	�9.+�9�T�9Xt�9��9͹�9���9��9���9���9���9���9#��9a��9���9x   x   v��9Ǣ�9:g�9c/�9���9���9���9��9͆�9��9��9y��9(��9D��9+/�9�i�9���90��9��9U�9��9��9O��9Q��9u��9���9Х�9΃�9�U�9��9x   x   �"�9U��9���9�.�91��9���9^��9�j�9�[�9Xj�9���99��9��98/�9��9���9%�9;|�9P��9��9bS�9��9���9���9B��9��9�R�9��9���9�{�9x   x   g8�9)��9}i�9>
�9ĺ�9l}�9�I�9�5�9�6�9�G�9�|�90��9f	�9�i�9���9�8�9ܭ�99�93x�9���9��9�D�9�T�90V�9�B�9��9���9�x�9��9���9x   x   �$�9��9�*�9���9j�9r(�9x��9E��9x��9c)�9�j�9ݽ�9Q+�9��9%�9��9h*�9+��9��9�u�9K��91��9G��9N��9=��9�t�9��9Ԫ�9~)�9���9x   x   ���9�U�9��9=S�9L��9���9w��9���9?��9>��9jS�9��9�T�9Q��9X|�9I�98��9G8�9��9��9^F�9�g�9�g�9�E�9�9+��9�9�9߬�9��9 |�9x   x   �r�9���92P�9���9���9�O�9@D�9�P�9��9+��9JO�9v��9�t�9��9u��9Lx�9��9��9� �90}�9$��9���9J��9�{�9"�97��9H�9'y�9w��9�9x   x   ���9::�9���9�B�9��9B��9p��9u��9�B�9���9�:�9f��9?��9>U�9��9���9�u�9��9@}�9���9m��9���9��9B~�9��97x�9/��9��9T�9_��9x   x   �.�9���9K�9w��9�_�9+G�9*`�9ǜ�9*�9G��9�.�9;��9��9Ă�9�S�9��9s��9xF�9>��9s��9m�95��9��9�G�9��9;�9�R�9Ą�9���9���9x   x   ^h�9���9"I�9���9��9���9���9]I�9���9Xg�9v"�9���9.��9_��9'��9�D�9c��9�g�9���9���9>��9��9Kh�9B��9�C�9a��9ӥ�9R��9 ��9�!�9x   x   1��9] �9��9�C�9n/�9{E�9B��9� �9z��9�I�9��9���9e��9���9��9�T�9}��9*h�9t��9-��9��9Vh�9��9|V�9���9V��9���9���9��9�I�9x   x   ��9q3�99��9���9+��9���9�3�9.��9Ok�9U4�9�9�9���9���9��9tV�9���9�E�9�{�9Y~�9�G�9J��9|V�9��9T��9L��9;�9�9Z5�9�j�9x   x   ���9�p�9"�9V�9�"�9`q�9J��9Ƀ�9PM�9�(�9�9\�9;��9���9���9 C�9u��9?�9="�9	�9��9�C�9��9Z��9���94�9��9a(�9�L�9v��9x   x   &�9���9N��9v��9��9<$�9���9�i�9i;�9��9��9f�9���9E��9_��9��9�t�9Z��9]��9Tx�9M�9r��9]��9K��94�9��9��9�;�9/j�9��9x   x   �z�9�-�9(�9w,�9m}�9d��9���9�X�9C1�9��9A�9��9G��9*��92S�9���94�9�9�9j�9Q��9�R�9��9���94�9��9��9y2�9�W�9S��9���9x   x   ���9��9���9?��9fK�9D��9���9X�9}<�9d'�9��9Y��9t��9��9@�9�x�9��9��9Hy�9��9τ�9U��9���9�9[(�9�;�9�W�9 ��9��9L�9x   x   r{�9\`�9E|�9���92�9E��9n��9bi�9�M�9r4�90�9���9���9?V�9���9�9�)�9�9���93T�9���9��9��9N5�9�L�9"j�9H��9��9A1�9���9x   x   :�9^8�9�j�9���9.I�9���9���9���9&k�9�J�9�"�9|��9ҙ�9��9�{�9���9ޮ�9?|�9-�9k��9���9�!�9�I�9pj�9f��9
��9���9�K�9���9xi�9x   x   U0�9�B�9C��9��9=��9���9���9u��94��9���9،�9�g�9�9��9��9<�9���9��9	�9�f�97��9R��9���9��9ʎ�9!��9 ��9L�9��9�B�9x   x   �B�9�|�9T��9�i�9"$�9���9 ��9b��9��9#��9���9�X�9"��9�Z�9��9 ��9�Z�9���9IY�9���9_��9���9���9���9Q��9�$�9�l�9���9
|�9*@�9x   x   .��9D��9�M�9���9���9�s�9-T�9�8�9��9���9i��9�I�9;��92�9s�9��9���9H�9���9	��9u�9�9�9�U�9�t�9���95��9MK�9���9��9 �9x   x   k�9�i�9���9���9d2�9���9���9֠�94i�9'#�9���9{A�9���9x��9b��9Ę�9B�9M��9#�9j�9���9��9���9,3�9c��9X��9�l�9A�9D��9���9x   x   
��9 $�9���9V2�9~��9���9SU�9��9���9Y�9���93�9�p�9ֆ�9Dp�9p3�9���9�X�9B��9��9DW�9���9���9j1�9Q��9�!�9���9J��9�|�9��9x   x   ���9���9�s�9���9���9�7�9���9<z�9v�9ׅ�9��9�,�9kO�9;P�9.-�9D��9[��9�	�9$y�9���9�5�9z��9���9�s�9g��9���9BY�9�<�9�=�9kY�9x   x   o��9���9T�9���9:U�9���9^c�9���9X�9���9���9�$�956�9�#�9���9۱�9.V�9B��9�d�9���9�V�9���9�T�9���9���9HK�9<�9Q�9��9/L�9x   x   '��9/��9w8�9���9��9-z�9���9�I�9���9O��9#�9/�9 �9h�9���9X��9(J�9G��9ny�9��9R��9�8�9���9م�9�Q�9��9
�9�	�9��98R�9x   x   ��9���9W�9
i�9���9a�9X�9��9���9���9/�9m�9��9���9���9D��9�W�9Z	�9i��9i�9z�9_��9{��9�a�9{:�9( �9�92"�9>:�9a�9x   x   :��9���9���9�"�9�X�9ƅ�9~��9K��9���9D�9��9&�9+�9��9���9���9{��9JW�9`#�9���9"��9ؙ�9�{�9�[�9�H�96C�9�@�9H�9�\�9�|�9x   x   ���9C��9)��9���9i��9��9{��9�9-�9��9�!�9��9r�9��9���9��9���9=��9f��9"��9ō�9{��9�{�9p�92m�9kn�9�o�9�o�9cz�9߇�9x   x   �g�9kX�9RI�9IA�9�2�9�,�9�$�9%�9s�9.�9��9~�9!�9"#�9�+�9S3�9�A�9�G�9�Y�9f�9t�9,��9ċ�9���9W��9��9"��9��9<��9Kt�9x   x   ��9���9��9a��9�p�9[O�906�9
 �9��93�9|�9$�9�7�9�O�9�q�9ʗ�9��9��9��9H�9wc�9Ύ�9ȧ�9U��9��9���9��9[��9Yc�9*G�9x   x   ß�9�Z�9 �9[��9���9-P�9�#�9q�9��9��9��93#�9�O�9n��9w��9��9lZ�9Ϟ�9���932�9�e�9R��92��9���9e��9۳�9���9�g�93�9��9x   x   ���9���9J�9L��9>p�9/-�9���9���9��9��9���9,�9�q�9��9��9/��9J��9N]�9���9C�9�g�9���9���9+��9��9�9�g�9��9���9^]�9x   x    �9֌�9��9���9i3�9N��9��9s��9d��9��9<��9l3�9��9��98��9��9p��9� �9Y��9���9�L�9T��9��9+��98��9�K�9Y��9���9��9���9x   x   ���9lZ�9���9B�9���9n��9WV�9PJ�9%X�9���9���9�A�9(��9�Z�9d��9y��9�=�9��9.^�9f��9��9W�9�c�9V�9��9��9=\�9���9>�9<��9x   x   ٞ�9���9H�9_��9�X�9�	�9g��9v��9�	�9W�9��9H�99��9 ��9r]�9� �9��9�w�9�	�9�9��9���9N��9���9��9�
�9ox�9W��9P�9F]�9x   x   ��9AY�9���9##�9`��9Sy�9�d�9�y�9���9�#�9���9�Y�9�9���9���9���9C^�9�	�9���9��9�P�9�m�9#Q�9�9Ö�9
�9�[�9Ɣ�9���9��9x   x   �f�9��9��9'j�9��9-��9���9��9Ui�9���9r��9`f�9qH�9o2�9x�9���9���9+�9��9�i�9��9���9Dk�9��9�}�9���9T��9��9�0�9�I�9x   x   F��9r��9��9��9{W�9�5�9W�9���9��9���9��9kt�9�c�9Hf�9h�96M�9��9:��9�P�9��9���9ƞ�9�M�95��9��9\L�9�g�9�h�9�c�9�s�9x   x   f��9��9�9�9I��9ޞ�9Ý�9N��9�8�9���9A��9݇�9���9(��9���9
��9���9YW�9���9�m�9���9Ҟ�9�o�9e��9�W�9���9$��9���9���9��9���9x   x   ���9���9�U�9$��9@��9!��9U�9��9��9=|�9Z|�92��90��9���9��9N��9#d�9���9LQ�9^k�9�M�9o��9�b�9���9b��94��91��93��9|�9�|�9x   x   ���9���9�t�9j3�9�1�9�s�9$��9<��9b�9\�9�p�9f��9���9#��9���9}��9eV�9���9E�9��9M��9�W�9���9���9���9ܮ�9a��9�o�9�\�9 a�9x   x   ��9���9̣�9���9���9���9_��9R�9�:�9eI�9�m�9ʒ�9���9���9z��9���9)�9P��9��9(~�9�9���9n��9���9���9Ȓ�9o�9�I�9�:�9(R�9x   x   @��9�$�9u��9���9
"�9��9�K�9!�9� �9�C�9�n�9���9,��9C��9��9�K�9]��9�9>
�9���9xL�9,��96��9��9Ӓ�95n�9JB�9 �9P�9�I�9x   x   ��9�l�9}K�9m�9���9�Y�9��9l
�9v�9"A�9Wp�9���9V��9]��9�g�9���9�\�9�x�9�[�9}��9�g�9ǡ�9=��9`��9o�9FB�9k�9i	�9��9>Z�9x   x   e�9���9���9z�9���9�<�9��9�	�9�"�9�H�9p�9U��9č�9(h�9?�9���91��9���9��9��9�h�9���99��9�o�9�I�9 �9k	�9�9=�9i��9x   x   /��9,|�9��9w��9�|�9%>�9W�9��9�:�9�\�9�z�9���9�c�9o3�9B��9*�9M>�9��9���9�0�9�c�9��9|�9�\�9�:�9>�9��9=�9b{�9���9x   x   �B�9?@�9�9$��9T��9�Y�9zL�9�R�9ga�9*}�98��9�t�9�G�9g��9�]�9��9m��9i]�9>��9�I�9�s�9���9�|�9a�9R�9�I�9/Z�9`��9���9�~�9x   x   d��9h�9�i�9
�90��9��9��9YE�9��9��9=��9���9���9�x�9���9C �9���9 x�9d��9���9���9Ծ�9��9�E�9��9k��9���9t	�9]h�9F�9x   x   Z�9"A�9��9o�9�Q�9LS�9�p�9���9��9a��9,�9���90��9-�9�Z�9lZ�9 �9��9���9��9��9h��9��9q�9�P�9*Q�9q�9���9�B�9�9x   x   �i�9ڻ�9K�9���9���9���9)��9��9+�9�+�9�9���9�d�9���9k��9��9nd�9���9,�9�*�9�+�9�9���9*��9w��9(��9�H�9ݺ�9j�9wJ�9x   x   �	�9�n�9���9a��9���9��9���9��9ۇ�9vi�9�4�9��9$4�9�n�9�o�9d4�9���94�9j�9%��9���9���9��9)��9<��9���9Rr�9��9���9e��9x   x   ���9�Q�9���9���9]l�9�G�9�/�9�9���9A��9!B�98��9��9?�97�9���9=B�9Χ�9:��9$�9�0�9�H�9�l�9���9���9�N�9	��96��9��9���9x   x   ���9S�9���9��9�G�9F�9���9��9O�9S��9�Z�9���9���9���9��9�Z�9���9�O�9
��9���9#�9�G�9ۏ�9��9#S�9���9a��9�d�9�f�9��9x   x   m�9Dp�9���9���9s/�9���9���9��9+��9K �9�w�9���9���9���9�v�9:!�91��9^�9��9��9	1�9|��9���9�n�9��9���9���9ks�9M��9��9x   x   �D�9���9��9���9`�9՚�9��9ǌ�9Y��9�M�9*��9���9ũ�9��9M�9���9ь�9��9w��9<�9���9��9B��9�D�9J��9���9���9���9̽�9��9x   x   ���9���9�*�9���9���9�N�9��9N��9�@�9[w�9���9���9'��93x�9@�9;��9ԫ�9�O�9��9
��9�,�9��9d��9�F�9A�9���9���9���9]�9uF�9x   x   ���9	��9�+�9Ai�9��90��9. �9�M�9Vw�9���9Ɵ�9B��9C��9�w�9N�9� �9_��9���9j�9)�9���9L��9ޔ�9�r�9�]�9�N�9�J�9^�9$u�9���9x   x   ���9� �9��9�4�9�A�9zZ�9�w�9)��9���9ğ�9���9ʟ�9���9��9�v�9"[�9XC�9G4�9��9< �9���9?��9S��91��93��9���9���9k��9���9���9x   x   "��97��9���9���9��9���9���9��9���9=��9ß�9(��9��9`��9m��9���9��9��9���9/��9��9��9��9t*�9�-�9�-�9\)�9��9��9��9x   x   B��9ݙ�9�d�9�3�9��9���9���9ǩ�92��9Q��9���9��9*��9���9�9�3�9�f�9���9���9Z �9o9�9<^�9&v�9ˑ�9Q��9��9w�9�[�9�8�9# �9x   x   ]x�9��9���9�n�9�9���9��9$��9Cx�9�w�9���9k��9���9��9o�9���9m�9�y�9U��9�$�9�n�9���9��9���9��9\��9���9:q�9r%�9���9x   x   D��9wZ�9C��9�o�9&�9��9�v�9)M�9)@�95N�9�v�9���9/�9#o�9#��9Z�9F��9�]�9f��9mE�9?��9���9c�9��9`�9��9��9�B�9_��9�^�9x   x    �9BZ�9��9W4�9���9�Z�9L!�9��9f��9� �9O[�9���9�3�9���92Z�9=�9��9�E�9���9t]�93��9��9-�9-�9n�9���9�^�9���9�C�9��9x   x   s��9��9^d�9���9BB�9���9Q��9��9��9���9�C�96��9�f�9��9Z��9���9`i�9�(�9d��9y\�9B��9��9^�9��9���9v[�9,��9�(�9�j�9��9x   x   �w�9��9���9'4�9��9P�9��90�9AP�9:��9�4�9U��9��9	z�9�]�9�E�9�(�9���9ǫ�9(7�9��9 ��9���9���9�8�9׬�9���9�(�9�C�9t^�9x   x   Q��9���9<�95j�9e��9=��9E��9���9c��9Wj�9=�9��9F��9���9���9 ��9~��9ګ�99c�9N��9_<�9Q�9�:�9t��9+a�9��9���98��9���9���9x   x   ���9��9�*�9Q��9V�9��9f��9��9j��9�)�9� �9���9� �9L%�9�E�9�]�9�\�9L7�9Y��9�`�9���9���9]b�9���9�7�9#]�9�]�9�D�9�#�9��9x   x   ���9%��9�+�9֑�91�9t�9g1�9C��9V-�9@��9��9:�9�9�9*o�9���9���9{��9��9z<�9���9J��9U��9�9�9���9/��9y��9t��9�q�9s:�9��9x   x   ��9���9,�9���9I�9�G�9��9��9���9���9���9j�9�^�9���91��9�9��9\��9:Q�9Р�9^��9#S�9S��9��9�9���9���9J\�9S�9u��9x   x   ,��9:��9���9'��9m�9>��9I��9���9߄�9]��9���9+�9�v�9w��9��9u-�9��9���9;�9�b�9�9�9_��9x�9�-�9��9;��9�x�9V�9���9���9x   x   �E�9�q�9l��9x��9��9���9]o�9/E�9G�9ss�9���9�*�9X��9Z��9G�9l-�9��9��9���9���9���9��9�-�9q�9���9���9�)�9���9t�9�F�9x   x   ��9Q�9���9���94��9�S�9�9���9��9G^�9���9N.�9Օ�9���9��9��9>��949�9ca�9 8�9Q��9%�9��9���9z��9�/�9���9�_�9n�9���9x   x   ���9]Q�9e��9���9�N�9��92��9��9!��9O�9��9^.�9���9���9���9��9�[�9-��9X��9J]�9���9���9J��9���9�/�9Ҿ�9�M�9I��9���9���9x   x   ��9Hq�9�H�9�r�9e��9ˎ�94��9��9r��9�K�9��9�)�9�w�9��9b��90_�9}��9���9��9�]�9���9���9�x�9�)�9���9�M�9��9���9��9��9x   x   �	�9ּ�9!��9��9���9�d�9�s�9��9q��9�^�9���9'�9O\�9�q�9C�9���9)�9�(�9o��9�D�9�q�9P\�9X�9���9�_�9=��9���95u�9�f�9��9x   x   sh�9�B�9Aj�9:��9Z��9%g�9���9C��9��9�u�9Y��9z�9S9�9�%�9���9�C�9=k�9?D�9���9�#�9�:�9Z�9���9t�9Z�9���9��9zf�9+�9���9x   x   T�92�9�J�9���9?��91��9H��9z��9�F�9+��9��9!�9� �9���9�^�9/��91��9�^�9���9��9��9n��9���9�F�9���9w��9��9ϖ�9���9�J�9x   x   S=�9�n�9���9Ӧ�9˩�9%��9�F�9&��9 [�9���9oI�9��9��9�f�9e��9c�9���9�f�9M��9 ��9!J�9k��9�[�9���9jG�9���9̨�9��9���9�n�9x   x   �n�9���9�I�98�9s.�9�u�9���9�B�9D��9@�9�[�9�{�9�^�9���9vB�9�C�9���9�]�9�{�9�Z�9)�9v��9�@�9^��9�s�9X-�9W�9�J�9)��9"o�9x   x   ���9�I�9��9���9"��9K"�9{q�9��9� �9d�9�~�9&g�9��9���9���9[��9B�9h�9i�9`c�9��9���9dq�9�!�9���9x��9��9�H�9f��9z��9x   x   ���9�9���9���9���9L��9�2�9Jj�9���9���9��9S�96��9Y�9��9{��9~S�9%��9;��9��9ii�9a3�9���9���9���9���9� �9��9(g�9�d�9x   x   ���9>.�9��9y��9z��9[��9'��9
�9F�9���9ӻ�9{P�9��9þ�9c��9�N�9���9��9�9{
�9���9���9��9���9Y��9�+�9���9(V�9<�9|V�9x   x   ���9xu�9"�9)��9C��9���9���9'��9��9[C�9���9z=�9 y�94x�9?�9E��9�A�9���9��9���9��9���9o��9�!�9�t�9H��9���9�M�9�O�9V��9x   x   eF�9���9Aq�9�2�9��9���9}��9R�9���9��9���9�4�9�G�9�4�9���9���9���9R�9��9���9&��9+3�9r�9���9DG�9��9���9���9���9���9x   x   ���9)B�9���9	j�9�	�9��9R�9~��9j�9~��98�9�+�9�+�9W�9���9�j�9:��9�R�9��9%	�9j�9���9IC�9'��9g�9�-�9E�9��9w-�9~g�9x   x   �Z�9��94 �9=��9�9؉�9���9j�9���9;��9��9k%�9��9p��9��9�i�9���9x��9��9���9� �9@��9�Y�9K�9x��9���9���9"��9!��9��9x   x   ��9��9�c�9H��9���97C�9���9x��93��9��9+�93,�9��9��9���9���9�A�9N��9��9Qb�9E�9I��90��9�}�9Pb�9�[�9Y�9�c�9��9��9x   x   �H�9)[�9�~�9���9���9|��9���9+�9��9+�9p7�98+�9S �95�9
��9P��9��9���9j�9MZ�9�G�95�9R)�9M�9��9��9��9�9�(�9D5�9x   x   ���90{�9�f�9�R�9JP�9[=�9�4�9�+�9j%�9A,�9@+�9%�9u+�9(7�9�=�9�M�9�R�9Uf�9J|�9���9G��9B��9���9���9���9��9���9@��9���9��9x   x   s��9t^�9p�9���9���9�x�9�G�9�+�9��9��9Y �9u+�9F�9x�9���9(��9��9�\�9S��9/��9��9aG�9Wk�9o��9���9���9!l�9;D�9E�9O��9x   x   �f�9���9`��9.�9���9)x�9�4�9e�9y��9��9R�9A7�9)x�9-��9^�9���9���9sh�9D��9�:�97��9���9z�9�'�9)�9!�9���9=��9�9�9���9x   x    ��9(B�9c��9��9P��9?�9���9���9��9���9/��9�=�9��9c�9L��9�B�9���9��9��9���9��9�_�9��9���93��9�]�9*�9ȟ�9
�9:��9x   x   �9�C�93��9g��9�N�9W��9���9�j�9�i�9̉�9��9�M�9Q��9���9�B�9��9h��9l��9^X�9���9�r�9��9��9%��9���9t�9_��9�Y�9:��9��9x   x   o��9���9,�9|S�9ż�9B�9���9y��9���9�A�9e��9%S�9��9 ��9��9���9��9���9��9>'�9k��9T��9	!�9P��9 ��9='�9K�9K��9/��9���9x   x   �f�9�]�9h�9/��94��9Ê�9NR�9S�9Ŋ�9���9��9�f�9]�9�h�9D��9���9���9=��9���9�:�9x��9���9���9���9�;�9���9���9��9���9���9x   x   6��9�{�9w�9T��9G�9T��9`��9`��9O�9W��9��9�|�9���9���9�9�X�9��9���9`o�96�9���9V��9~�9m�9�m�9w��9���9�Y�9��9n��9x   x   ��9[�9~c�9��9�
�9=��9��9�	�9��9�b�9�Z�9��9���9>;�9Y��9���9p'�9�:�9H�9���9*��9x��9���9\�9�<�9�&�9���9ݠ�9[9�9i��9x   x   -J�9C�9��9�i�9%��9d��9���9�j�9n!�9��9-H�9Ч�9Q�9���9�9%s�9���9���9ـ�95��9�9��9��9z��9���9�s�9��9×�9��9��9x   x   ���9���9��9�3�9��9h��9�3�9��9Ұ�9���9�5�9Դ�9�G�9��9M`�9���9���9<��9���9���9%��9��9n��9���9���9<`�9B��9jE�9D��9�6�9x   x   �[�9�@�9�q�9���9p��9���9�r�9�C�9bZ�9Ӫ�9�)�9&��9�k�9�9l��9|��9i!�97��9Y~�9Ϭ�9��9���9j �9v��9���99�9{m�9f��9�)�9���9x   x   !��9���99"�9 ��9Q��9("�9"��9���9��9�~�9��9X��9��9>(�9)��9���9���9��9��9��9���9���9���9��9P)�9���9���9��9�~�9\�9x   x   �G�9�s�9��9=��9���9.u�9�G�9�g�9��9�b�9��9���9[��9�)�9ș�9,��9n��9J<�9 n�9�<�9���9���9���9T)�9w��9=��9�9�d�9���9de�9x   x   ���9�-�9���9���9R,�9���9���9�.�9N��9�\�9C�9���9>��9��9\^�9�t�9�'�9]��9�9'�9t�9Y`�9L�9���9:��9��9�[�9í�9>1�9 ��9x   x   ���9��9X��9� �9&��90��9$��9��9C��9�Y�9��9@��9�l�9��9��9���9��9���9Ѐ�9���9��9W��9�m�9���9��9�[�9m��9&�9[��9�9x   x   ��9�J�9.I�9n��9�V�92N�9��9n�9±�9�d�9��9���9�D�9ϗ�9P��9Z�9���9ϵ�9�Y�9��9ݗ�9wE�9l��9��9�d�9���9�9���94P�9�V�9x   x   ��9M��9���9vg�9`<�9+P�9s��9 .�9���9{��97)�9 ��9��98:�9��9���9���9��9�9}9�9��9G��9y)�9�~�9���9'1�9E��90P�9t:�92g�9x   x   �n�9Bo�9���9!e�9�V�9���9T��9�g�9:�9���9�5�9~��9���9��9���9w��9E��9���9���9��9��9�6�9u��9=�9Ke�9���9���9�V�9$g�9���9x   x   g4�9e�9���9���9��93��9TT�90(�9w�9_��9/��9�4�9�|�9Jt�9��9�E�9��9�t�9�}�9�5�9���9;��9��9�)�9�T�9��9z�9Z��9���9�d�9x   x    e�9��9�y�9#{�9���9yN�9���9���9��9\6�98��9��9_+�94��9�N�9eP�9��9%*�9��9���9�8�9��9`��9���9N�9���9:{�9�z�9R��9[e�9x   x   ���9~y�9y?�9U�9[��9'�9���9�h�9�9���96��9�9��9�e�9���9�c�9l��9$�9M��9ӊ�9�9�h�9,��9h&�9��9�U�9>�9Py�9-��9��9x   x   ���9�z�9�T�9�m�9m��9�"�9���9��95��9t��9��9\��9��9���9��9z��9���9��9���9ǎ�9��9ǟ�9K"�9 ��9Gl�9V�9y{�9M��9?��9��9x   x   ��9���9'��9U��9���9�<�9t��9'��9�)�9!J�9�5�9���9XQ�9xy�9�P�9���9�6�9�K�9�'�9Q��9���9h<�9G��9���9y��9,��9��9b��9���9ö�9x   x   ˚�9+N�9�&�9�"�9�<�9rd�9��9յ�9��9���9wX�9���9�9&�9���9LY�9
��9���9��9=��9"f�9N=�9\!�9�'�9EM�9���9X'�9q��9���9�%�9x   x   �S�9c��9���9���9M��9��95��99w�90E�9��9p}�91��9���9���9+|�9e��9lE�9�v�9��9x��9Ɨ�9m��9��9&��9�T�9���9ގ�9Gx�9���9���9x   x   �'�9��9-h�9e�9���9���9+w�9�,�9���9eB�9Ɲ�9���9���9\��9�B�9���9�,�9	w�9��9���9  �9�g�9���9�'�9���9
h�9�@�9�A�9Yg�9���9x   x   ��9���9��9��9�)�9���9E�9���9k3�9���9ݷ�9���9̷�9���9�1�9 ��9=F�9ֽ�9y(�9���9��9Q��9��9X��9"i�9!8�9"0�98�9�h�9���9x   x   ���9�5�9���9&��9�I�9Ȧ�9���9WB�9���9���9���9��9o��9<��9$E�9q��9��9AK�9���9���9�7�9T��9`��9�x�9Q�9�A�9�@�9�R�9\x�9i��9x   x   ���9���9���9��9�5�9CX�9S}�9���9Է�9���9���9��92��9f��9{�9jZ�9�5�9e�9r��9/��9���9m��9|y�9�k�9�e�9�d�99e�9bj�93z�9T��9x   x   `4�9t�9��9	��9d��9^��9#��9���9���9���9��9!��9���9,��9���9���9f��9�9�9w4�9rK�9�_�9�s�9��9���9Ō�9\��9�t�9�_�9#I�9x   x   c|�9�*�9���9���9'Q�9�9q��9���9ҷ�9|��9?��9���9���9�9�P�9D��9���9�)�96}�9`��9�	�9RP�9d��9���9��9'��9b��9�M�9T�9���9x   x   �s�9���9�e�9U��9Oy�9�9���9f��9��9`��9���9?��9�94z�99��9?d�9M��9�s�9w �9�}�9���9�J�9z�9ɝ�9���9�z�9$L�9���97{�9J �9x   x   �9+N�9@��9V��9�P�9���9;|�9�B�9�1�9NE�9.{�9��9Q�9K��9���9O�9��9O��9���9�,�9S��9�$�9�c�9�~�9�c�9�"�9g��9�,�90��9���9x   x   lE�9P�9nc�9c��9���9SY�9���9���9:��9���9�Z�9���9u��9cd�9)O�9�D�9;�93�9��9��9Pm�9���9��9��9���9�m�9��9L�9C1�9=9�9x   x   ��9���9Q��9���97�91��9�E�9�,�9�F�9l��96�9���9���9���9��90;�9sg�9���9<��9 Z�9���9"U�9�v�9�T�9x��9[�9��9���9@k�9);�9x   x   wt�9*�9&�9��9L�9���9�v�9`w�9:��9�K�9��9{�9*�9Ft�9���9<3�9���93��9���9���9�:�9���9Ɇ�9;�9���91��9���9H��9h0�9���9x   x   �}�9��9a��9���9�'�9j��9]��9`��9�(�9��9���9��9�}�9� �9��9��9e��9���9���9���9�-�9i[�9P,�9���9J��9���9ц�9C�9I��9 �9x   x   |5�9���9���9��9���9���9��9��9���9���9���95�9���9�~�9�,�9o��9lZ�9��9ϳ�9�d�9k��9N��9�d�9���9��9�Y�9���9�,�9�|�9���9x   x   Ǩ�9�8�9R�9 �9��9�f�9Q��9� �96�9_8�9!��9L�9s
�9H��9Ѿ�9�m�97��9�:�9�-�9|��9(�9���9�.�9:�9���99o�9���9���9?�9�J�9x   x   \��9?��9-i�9#��9�<�9�=�9��9�h�9��9��9��9R`�9 Q�95K�9S%�9��9�U�9��9�[�9x��9���9�Z�9���9�V�94��98$�9�K�9�O�9J_�9���9x   x   ��9���9}��9�"�9���9�!�9���9N��9Z�9'��9@z�9�t�9$��9�z�9qd�90�9Ew�9)��9�,�9e�9/�9���9
v�9�9xd�9M{�9��9xu�9�{�9˨�9x   x   �)�9>��9�&�9s��95��9-(�9���9T(�9!��9�y�9�l�9���9F��9���9��9f�9U�9�;�9	��9ܲ�9,:�9�V�9�9G�9��9G��9���9Vk�9x�9X��9x   x    U�9eN�9{��9�l�9��9�M�9�U�9���9�i�9�Q�9�f�9y��9Ш�9e��9Cd�9'��9	��9$��9���9I��9��9U��9�d�9��9���9q��9Tf�9�S�9�j�9��9x   x   Q��9$��9�U�9�V�9���9&��9���9�h�9�8�9�B�9�e�9���9��9S{�9k#�9�n�9�[�9���9���97Z�9no�9R$�9T{�9O��9r��9�d�9�B�9�6�9�i�9���9x   x   ��9�{�9y>�9�{�9u�9�'�9���9�A�9�0�9�A�9f�9*��9-��9�L�9��9���9���9���90��9���9۾�9�K�9��9���9Rf�9�B�9�1�9DB�9э�9G'�9x   x   ���9�z�9�y�9���9��9��9�x�9WB�9�8�9�S�9(k�9�u�9�N�9���9�-�9��9��9���9��9�,�9���9�O�9vu�9Ok�9�S�9�6�9DB�9|y�9���9Ķ�9x   x   ���9���9{��9���9��9��9G��9h�9Ai�9y�9�z�9�`�9	�9�{�9Ȋ�9�1�9�k�9�0�9���9}�9T�9O_�9�{�9x�9�j�9�i�9���9���9?��9��9x   x    e�9�e�9F��9Ӑ�9'��9h&�9h��9��9G��9��9��9�I�9���9� �9X��9�9�9�;�97��9E �9���9�J�9���9���99��9���9���9 '�9���9֑�9���9x   x   ]��9Z��9ƃ�9���9�'�9���9�
�9]I�9:��9/��9~��9+��9�}�9W��9�l�9C��9�i�9���9�~�9T��9���9���9Ú�9"K�9�
�9���9(�9'��9߃�9b��9x   x   <��9:A�9��9jb�9��9I��9���9���9�&�9�7�9�%�9���9V�9� �99y�9�z�9��9
�9F��9�$�9{9�9<(�9B��9t��99��95��9Ka�9��9l@�9���9x   x   ���9z�9��90l�9��9���9W��9���9��9��9:K�9��9���9X^�9֖�9]]�9���9��9�K�9��97��9���9��9���9��9l�9o�9
 �9���9�V�9x   x   u��9/b�9l�9+��9X�9��9Z��9��9r��9b�94��9��9�a�9���9r��9�b�9���9Q��9\�9��9o��98��9��9Y�9H��9�l�9B`�9��9`J�9]J�9x   x   A'�9���9P�9�W�9��97i�9�9��9P1�9g��9���9Љ�9��9�<�9a�9��9���94��9s/�9���9~�9`h�9���9�W�9k�9=��9P(�9��9�x�9��9x   x   "��9���9J��9^�9&i�9��9XD�9���9���9��9���9߄�92��9&��9s��9���9� �9���9��9�B�9���9j�9��9���9���9���9ym�9��9)�9lm�9x   x   N
�9S��9���9��9R�9@D�9gy�9���9��9*v�9<�9�w�9��9?x�9]�9^v�9Ġ�9՚�9�y�9%D�9)
�9S��9v��9���9e
�9�u�9��9���9\�9!u�9x   x   �H�9���9A��9���9Ю�9g��9���9v�9�1�9���9i3�97q�92q�93�9���9�1�9�u�9���9��9D��9e��9��9���9�H�9���9]�9�3�94�9�\�9���9x   x   ���9'&�9���9��91�9w��9���9r1�9l��9Q �9�V�9�q�9]V�9w!�9���9q0�9��9��9�.�9��9���9i'�9���9�#�9c��9���9b��9J��9���9�$�9x   x   x��9�6�9���9��9��9j�9v�9p��9V �9VX�9�k�9dl�9lW�9��9���9�t�9(�9���9a�9ۦ�9�7�9���9Î�9�P�94,�9��9��9�,�9�N�9{��9x   x   ���9%�9�J�9ɂ�9���9���9�9W3�9�V�9�k�9]i�9l�9	X�92�9>�9{��9���9f��9ZI�9Q%�9r��9��9���9%��9��9���9۶�9���9d��9���9x   x   x��9���9p��9���9���9���9�w�9'q�9�q�9el�9l�9Xp�9Nq�9nx�9ӄ�92��9>��9��93��9���9(�9H'�93�9�G�9�L�9M�9H�9k2�9�&�9� �9x   x   $}�9��9��9\a�9��9��9��94q�9vV�9uW�9X�9eq�9���9d��9��9�b�9���9"�9�~�9���9h8�9)|�9���9���9%��9���9ϳ�9|�9�:�9��9x   x   ���9J �9�]�9r��9�<�9��9Cx�93�9�!�9��9-2�9�x�9m��9a>�9���9`^�9��9��9L�9~��9}r�9��98-�9^U�9\U�9-�9���9q�9���9�L�9x   x   Ml�9�x�9���9A��9G�9s��9w�9���9���9��9t�9��9��9���9��9=y�9Zk�9�T�9`6�9��9R��9�/�9d��9���9Հ�9/�92��9R�9�6�95T�9x   x   ͤ�9�z�9$]�9zb�9#��9��9�v�92�9�0�9�t�9���9y��9�b�9�^�9Sy�91��9S��9f�9��9��9��9T�9ړ�9.��90T�9���9~�9��9��9���9x   x   �i�9��9׸�9���9ͨ�9�9��9Cv�9l��9��9���9���9ж�9�9�k�9h��9�N�9=��9���9m��9Ƨ�9�(�9�O�9H)�9��9k��9 ��9��9Q�9w��9x   x   W��9��9��9]��9a��9*��93��9��9���9��9ށ�9���9��9e��9U�9��9V��9�'�9�w�9�|�99�9_��9���9R8�9�{�9�v�9`)�9���9l�9�U�9x   x   �~�9A��9L�9��9�/�9~��9}z�9���9�/�9 �9�I�9���9Y�9�L�9�6�9K�9���9�w�9��9��9i�9J��9�i�9��9���9	v�9K��9��9[7�9iK�9x   x   W��9%�9��91��9
��92C�9�D�9ް�9���9���9&�9a��9N��9��9g�9I�9���9�|�9"��9���9-#�9�"�9j��9~��9�~�9��92�9?�9���9��9x   x   ���9�9�9}��9׶�9��9(��9�
�9$��9l��9�8�9B��9��9,9�9/s�9��9���9+��9e9�9>i�9F#�9�j�9�#�9�k�98�9���9���9%��9Mq�9:�95�9x   x   ��9{(�9A��9���9�h�9#k�9��9���9:(�9���9 ��9&(�9�|�9���9P0�9�T�9<)�9ɞ�9���9,#�9�#�9_��9Ǟ�9f+�9�S�9!.�9P��9�}�9�&�9���9x   x   ���9���9m��9L�90��9X�9@��9���9���9���9���9 4�9���9.�9.��9���9vP�9q��9-j�9���9�k�9מ�9�N�9Y��9���9{-�9s��9�3�9��9F��9x   x   ^K�9���9n��9�Y�9�X�9n��9i��9zI�9�$�9�Q�9%��9�H�9���9FV�9���9��9�)�9�8�9���9���9H8�9+�9^��9Ē�9&V�9���9I�9K��9�O�9%�9x   x   �
�9���9��9���9�9���9>�9p��9[��9:-�9���9�M�9��9JV�9���9�T�9���9{|�9Y��9�9��9�S�9���9,V�9���9nM�94��9�-�9���9��9x   x   6��9���9�l�9m�9���9���9[v�9^�9���9��9���9N�9���9.�9�/�9m��9��9ow�9�v�9]��9���9L.�9�-�9���9nM�9b��9��9���9Y]�9w�9x   x   W(�9�a�9��9�`�9�(�9<n�9h�9m4�9T��9��9��9I�9Ǵ�9w��9��9?�9���9�)�9���9��9`��9t��9���9!I�95��9��9���9�4�9!�9#n�9x   x   c��9' �9u �9j��9���9r�9���9�4�95��9�-�9���9Z3�9�|�9�q�9�9��9~��9���9U�9��9wq�9�}�9�3�9G��9�-�9���9�4�9`��9R�9z��9x   x   ��9�@�9��9�J�9{y�9��9�9�]�9���9�O�9N��9m'�9�;�9���9S7�9]	�9�Q�9��9�7�9���9:�9�&�9��9�O�9���9?]�9�9@�9�y�9DJ�9x   x   m��9���9�V�9�J�9���9n�9�u�9y��9�%�9G��9\��9��9���9�M�9�T�9��9���9�U�9�K�9*��9@�9���9&��9�$�9ۻ�9�v�9�m�9T��96J�9qW�9x   x   �Q�9���9=x�9���9��9-��9~p�9�#�9|��9p��9N\�9D��9Л�9X�9���9�E�9���9i�9���9ݫ�9\�9n��9��9�%�9�n�9���9���9���9�z�9���9x   x   ���9�2�9�6�9r��9Y��9m��94d�9j��9��9�.�9s��9=��9�&�9c>�9���9a��9�>�9�$�9��9��9�.�97��9��9�b�9���9p��9���9}5�9�0�9ϣ�9x   x   x�9�6�9�f�9� �9���9�%�9F��9��9�f�9���9F��9}i�9��9��9q��9��9��9�j�9��9��9kf�97��9���9�%�9���9 �9�i�9�7�98x�9�5�9x   x   |��94��9� �9���9���9H��9���9�9�D�9]A�9���9�Q�9�A�9��9Ϻ�9�A�9$R�9���9�A�9�E�9�9���9��9���9��9���9���9~��9�`�9&b�9x   x   t��9���9D��9{��9�K�9~I�9nK�9IF�9�*�9���9�?�98J�9���9�"�9���97I�9@�9R��9�)�9_E�9�L�9�H�9�J�9���9���9Ɲ�9���9��9���9�9x   x   ���9���9{%�9���9`I�9y�9���9�{�9
�9e�9�x�9�2�9̟�9���9T2�9�y�9�c�9a�9�}�9H��9��9J�9���9[&�9���9���92�9���98��9�3�9x   x   �o�9�c�9Ո�99��9;K�9���9�A�9���9`��92��9���9�,�9�]�9�-�9?��9���9���9���96A�9]��9�J�9���9���9d�9n�9?��9�D�9��9�E�9Q��9x   x   0#�9���9���9��9�E�9k{�9���9��9ͩ�9_c�9���9�.�9y.�9���9^c�9s��9и�9Y��9�|�9�F�9~�9b��9L��9L$�9�u�9�
�9z��9o��9��9�u�9x   x   ���9Y��9f�97D�9�*�9��9B��9ũ�9=K�9k��96�9�)�9#�9��9�K�9٨�9���9�
�9�(�9~D�9oe�95��9���9�f�9���9ο�9���9��9��9�f�9x   x   ���9�-�9#��9�@�9���9�d�9��9Hc�9d��9I�9w1�9�1�9��9 ��9�d�9D��9 d�9���9^A�9���9�,�9ֽ�9�Y�9�9���9���91��9��93�9�Y�9x   x   b[�9���9���9v��9q?�9[x�9[��9���9-�9{1�9yD�9�1�9��9���9ˬ�9�y�9�>�9 ��9w��9���9�[�9�3�9y�9��9���93��9#��9��9(�9�2�9x   x   b��9��9�h�9uQ�9�I�9�2�9�,�9�.�9�)�9�1�9�1�9�'�9�.�9�-�9r2�9�I�9�Q�9Ek�9Ň�9:��9���9���9��9��9d*�9c*�9��9��9T��9���9x   x   ���9�%�9���9SA�9���9���9�]�9{.�95�9��9��9
/�9�\�9'��92��9B�99��9L%�9��9:�9�x�9T��9p�9^H�9�O�9�H�9q�9o��9�w�9s�9x   x   ��9�=�9��9Ȼ�9Y"�9���9�-�9���91��9K��9���9�-�9>��9�#�9���9��97?�9��9Z��9֑�9�@�9P��9
&�9�T�9(T�9�$�9���9 ?�9���9J��9x   x    ��9=��9��9���9^��9K2�9c��9�c�9�K�9,e�9��9�2�9]��9���9K��9g��9n��9�9�0�9�*�9F�9|��9���9�$�9���9��9+�9Q,�9�-�9��9x   x   dE�9���9��9�A�9=I�9�y�9��9ĩ�9.��9���9�y�9J�9�B�9N��9���9�F�9j��9�%�9��9"��9=��9�6�9���9���9�4�9ח�9���9{�9E)�9��9x   x   '��9�>�9��9!R�9)@�9�c�9&��9C��9 ��9xd�9?�9qR�9���9�?�9���9���9g}�9f.�9��9���9c��9�{�9ʯ�9~�9���9���9.��9x-�9(|�9-��9x   x   �9�$�9�j�9���9���9��93��9��9g�9l��9���9�k�9�%�9�9b�9#&�9�.�9�
�9Ǩ�9���9���9�K�9�I�9P��9+��9c��9&�9�-�9�&�9N�9x   x   ֜�9߈�93��9 B�9+*�9~�9�A�9n}�9)�9B�92��9~��9Λ�9���91�9s��9j��9��9�O�9��9'P�9��9gR�9���9�P�9o��9���9���9�.�9>��9x   x   ֫�98��9W��9�E�9�E�9���9��9�G�9QE�9���9���9��9�9���9W+�9���9���9��9-��9Y��9>5�9v4�9���9��9@��9K��9���9�+�9{��9'�9x   x   \�9�.�9�f�9��9&M�9��9�K�9a�9^f�9�-�9�\�9���9�y�9�A�9�9��9���9-��9jP�9\5�9�|�9�5�9AS�9���9$��9��9)�9>�9]x�9���9x   x   ���9���9���9c��95I�9�J�9���9W��9C��9��9 5�9���9f��9J��9\��9�7�9~|�9pL�9F��9�4�9�5�9��9�K�9�~�9�5�9���9���9���94��9�3�9x   x   `��9~��9���9���9SK�9���9���9\��9���9�Z�9��9��9��9'�9w��9q��9���9lJ�9�R�9��9qS�9�K�9N��9��9:�9�%�9j�9e�9$�9�\�9x   x   �%�9]c�9&�9H��9Ă�9H'�9e�9`%�9h�9=�9��9� �9�I�9�U�9�%�9���9�~�9���9.��9{��9���9#�9��9�#�9U�9]K�9!�9:�9�9�f�9x   x   �n�9C��9C��9͝�9���9���9!o�9�v�9���9"��9���9�+�9�P�9IU�9� �9�5�9^��9���9#Q�9���9p��9�5�9S�9U�9�P�9�*�9]��9N��9+ �9bw�9x   x   ���9��9� �9[ �9���9���9C��9��9��9���9q��9�+�9J�9	&�9��9˘�9���9��9���9���98��9,��9�%�9fK�9*�9��92��9S��9�
�9
��9x   x   G��9���9�j�9j��9���9	3�9�E�9���9ˡ�9j��9[��9� �9��9���9:�9��9���9��9(��9��9m�9��9|�9!�9Z��9*��9��95��9�F�9�3�9x   x   <��9�5�98�9��9��9���9� �9y��98��9B��9�9��9���9@�9L-�9Z��9=.�9�.�90��9L,�9K>�9���9r�9'�9@��9?��9��9 !�9��9�9x   x   �z�91�9�x�9ha�9���9��9�F�9��9  �9H�9@�9m��9�x�9���9�.�9*�9�|�9a'�9/�9���9�x�9@��9�9��9
 �9�
�9�F�9��9Y��9na�9x   x   ��9
��96�9�b�9��9|4�9��9sv�9�g�9�Z�9�3�9���9h�9.��9��9���9���9��9���9Q�9���9�3�9�\�9�f�9#w�9ҷ�9�3�9��9Wa�9�4�9x   x   �J�9p��9���95V�9���9�=�9�K�9���9�9!r�9���9��9���9$��9K��9&�9���9?��9���9��9K��9�r�9'�9���99I�9I;�9���9$V�90��9���9x   x   K��9VH�9`��9yf�9���9�n�9Px�9ҫ�9<��9��9]��9�X�94O�98��9�_�9�a�9\��99M�9�W�9u��9��9���9٭�9�w�9�q�9���9�d�9k��9F�99x   x   J��96��9���9���9$S�9?��9��9(��9���9���9|*�98�9���9޾�9x�9c��9E��9|:�9%*�9���9:��9���9-��9=��9�Q�9���9J��9Q��9^��9s]�9x   x   �U�9+f�9c��9���9FC�9u��9+��9"G�9���9�T�9Cq�9�9MG�9���9d��9�G�9)�9/p�9fU�9_��92F�9v��9���9�A�9L��9���9�b�9W�9`ý9JŽ9x   x   ��9$��9�R�9#C�9�y�9���9tI�9B��9��90�9��9�	�9k��9#�9���9l	�9���9��9S�9��9�J�9"��9�y�9�B�9�P�9-��9���9%ҿ9���9�ѿ9x   x   F=�9n�9���93��9���9��9��9�8�9p�9���9?�9���9�y�9�x�9b��9�9���9x�9l:�9� �9)��9��9z��9��9o�9�;�9�_�9���9$��9�a�9x   x   �J�9�w�9���9���92I�9��9��9��9c'�9v�9�i�9O��9�2�9� �9*j�9yu�9@)�9G��9���9 �9�K�9���9n��9�w�9�H�9�p�9���9���9���9�l�9x   x   ϡ�9���9���9�F�9��9�8�9���9���9��9��9��9���9���9��9	�9|�9+��9��9�9�9C��9�D�9���98��9���9u��9�D�9� �9|��9�F�97��9x   x   �9\��9���9n��9K�9/�9;'�9��9J��9a��9��9u �9_��9h��9���98�9�'�9��9�9��9j��9���9��9�h�9Z��9��9 ��9d��9:��9h�9x   x   q�9��9¦�9"T�9��9C��9Gv�9p�9\��9���9F��9f��9���9y��9	�9jv�9���9��9T�9���9}�9�r�9(��9��9d�9�E�9ZI�9�b�9���9���9x   x   t��9r��9�)�9�p�9���9��9�i�9���9��9O��9�9r��9~��95��9dh�9��9���9�o�9f)�9���9��9�y�9nU�9>�9j,�9G)�9'*�9�@�9�V�9�x�9x   x   �~�9�W�9�7�9z�9M	�9}��90��9���9p �9j��9x��9���9���9� �9k��9O�9K�9T9�9W�9;�9��9��9^��9��9�'�9�'�9��9��9���9���9x   x   ���9VN�98��9�F�9��9by�9�2�9��9r��9���9���9���9R1�9�x�9^��96H�9B��9{M�9���9Cv�9���9?b�9��9��9��9n��9��9g�9h��9}s�9x   x   9��9o��9I��9%��9��9�x�9� �9
��9���9���9i��9� �9�x�9��9���9���9t��9���9��9���9�Y�9�9.q�9���9��9�o�9���9:X�9x��9p��9x   x   |��9@_�9�9��9���9j��9Oj�9K	�9���9�	�9�h�9���9���9��9�9�_�93��9|(�9ց�9���9���9q~�9"��9�)�9���9��9���9��9@}�9�'�9x   x   ]%�9Pa�9��9�G�9q	�99�9�u�9��9��9�v�94�9��9�H�9��9�_�9^'�9���9e��9�Z�9���9���9X��9�'�9�&�9ƶ�9���9���9�Y�9��9g��9x   x   ��9��9��9�9���9&��9�)�9���9`(�9[��9���9��9���9߮�9y��9���9� �9�1�9�9���9���9���9��9N��9���9���9��9�1�9��9���9x   x   ��9M�9w:�9Vp�9*�9��9٤�9���9��9��9tp�9:�9,N�95��9�(�9���9�1�9�}�9�w�9��903�9i��9���9�1�9��9�w�9�}�9U1�9���9�(�9x   x   ���9�W�9K*�9�U�9��9;�9l��9�:�9��9U�9Q*�9�W�9k��9���9x��9%[�9g�9�w�9���9��9��9�T�96 �9��9��9(w�9��9L[�94~�9ؤ�9x   x   ��9���9��9���9���9@!�9��94��9���9���9���9A��9@w�9���9c��9���9~��9H�9��92l�9s#�9�"�9�i�9��9~�92��9���9���9���9�t�9x   x   b��9��9���9�F�9\K�9��9�L�9�E�9���9��9Q��9��9��9�Z�9���9n��93��9�3�9o��9�#�96��9$�9
 �9m2�9���9���9۵�9�V�9���9t��9x   x   �r�9��9���9+��9���9��9���9'��9���9t�9�z�9m��9~c�9C�9��9I��9���9��9$U�9#�9$$�9}S�9t��9r��9a��9 ~�9��9Jf�9��9Ny�9x   x   ��9I��9���9O��9�z�9���9���9|��94�9���9�V�9���9y��9|r�9Q��9�(�9���9���9� �9dj�9L �9���9}��9�'�9���9,q�9K��9G��9&U�9g��9x   x   !��9Ux�9���9�B�9�C�9(��9:y�9ݤ�9dj�9���9�?�9d�9v��9���9�*�9�'�9F��9�2�9{�9?�9�2�9���9�'�9�)�9���9��9I�9�B�9��9Yh�9x   x   �I�9pr�98R�9.��9�Q�9#p�9�I�9���9���9�e�9�-�9%)�9 
�9O��9��9��9���9q�9̓�9�9���9���9���9���9�9�'�9�+�9�c�9o��9���9x   x   �;�9��9}��9o��9.��9�<�9�q�9,F�9b��9RG�9�*�9J)�9���9\q�9]��9���9���9�x�9�w�9���92��9?~�9Pq�9)��9�'�9�-�9;H�9ϗ�9�D�9Lq�9x   x   ��9ne�9���9�c�9���9a�9���9��9���9�J�9�+�9M�9Y��9:�9״�9���9��9n~�9��9���99��9 �9]��9X�9�+�95H�9у�9�9���9Ib�9x   x   sV�9߇�9�9�W�9ӿ9���9.��9� �9ǔ�9Gd�9XB�9���9eh�9�Y�9P��9[�9�2�92�9�[�9^��9W�9rf�9H��9�B�9�c�9���9� �9n��9���9�п9x   x   i��9}F�9妼9Ľ9y��9��9���9�G�9���9J��9	X�9,��9���9���9^~�9Ӳ�9��9���9�~�9��9���9��9 U�9���9=��9�D�9u��9���9���9�Ľ9x   x   ੻91��9�]�9�Ž9@ҿ9�b�9�m�9Q��9Hi�9���9�y�9���9�t�9���9�(�9C��9c��96)�96��9�t�9}��95y�9=��9 h�9���9q�9b�9�п9aĽ9�[�9x   x   fN�9���9��9��9��9��9X��9x��9���9�	�9���9hm�9�S�9���95��9^Q�9��9��9�T�9an�9a��9
�9V��9���9K��9�9L��9��9���9���9x   x   U��9<��9�9
=�9R�9�a�91�9��9���9���9�9�9�@�9Ш�9�U�9�0�9�2�9^U�9���9q?�9�9�9��9���9���9R�9mc�9��9Z<�9�
�9P~�9׷�9x   x   g�9��9ɺ9�#�9��9�F�9���9>u�9�9���9���9��9���9((�9s��9�&�9��9��9���9���9��97t�97��9�F�9$�9"#�9˺9��9g��9���9x   x   �9�<�9r#�9���9
X�9��9���9�+�9lj�9b�9O��9��9�j�9�%�9�%�9�k�9��9m��9;b�9Lj�9�+�9���9���9.V�9牿9+"�9�:�9L�9�G�9vI�9x   x   Y��9��9?�9�W�9
�9��9L��9���9���9�G�9pV�9���9���9E4�9&��9���9X�9�G�9B��9���9w��9���9l�9�W�9��98�9렼9a��9�w�9"��9x   x   ��9�`�9F�9���9���9k��93�9��9<�9�'�92��9��9W|�9|�9���9^��9L'�9��9I��9�3�9q��9���9���9NF�9Ra�9��9@�9Rd�9�b�9��9x   x   K��9R�9��9 ��9���9�2�9�g�95��9�j�9��9e2�9���9u.�9t��9;3�9q �9�l�9���9|g�92�9���9l��9���9��9���9%��9^��9���9%��9��9x   x   K��9��9ut�9+�9@��9���9��9�.�9E��9|��9j|�9a��9���9�z�9̼�9���9h-�9܋�9��9���9�)�9�t�9���9���9<��9	�9ݯ�9o��9:�9ڶ�9x   x   ���9���92�9�i�98��9��9�j�91��9��9dZ�9>��9��9���9�Y�9n��9��9�k�9��9E��9.j�9��9��9L��9�9+n�9i�9)��9�9�n�9��9x   x   |�9e��9��9ea�9,G�9�'�9��9d��9dZ�9���9S�9��9]��9�Z�96��9��9�&�9�G�9`�9;��9���9��94y�9��94��9��9���9���9��9�y�9x   x   ���9e8�9���9���9�U�9���9*2�9I|�94��9_�9!�9m�9���9�{�9W1�9<��9�V�9|��9��9~8�9���9��9!��9�m�9�h�9jP�9�e�9go�9��9 ��9x   x   l�9�?�9��9E�9V��9���9���9Q��9��9��9}�9v�9���9y��9K��9x��9��9��9�>�99l�9��9��9���9Z�9�+�9,�9/!�9/��9���9ʞ�9x   x   �R�9ɧ�9���9j�9���9!|�9Y.�9���9���9z��9���9���9e.�9�{�9%��9�k�9Z��9��9KS�9���9��9U,�90��9A��9���9��9c��9�/�9f��9c��9x   x   ���9�T�9q'�9i%�9�3�9�{�9y��9�z�9Z�9�Z�9#|�9���9�{�9�4�9�$�9&�9�T�9���9���9���9`��9�9t5�9,�9�~�9K5�9ʛ�9���9���9���9x   x   6��9�/�9��9N%�9���9���9g3�9��9˜�9���9�1�9���9c��9�$�9���91�9���9E��9�:�9޻�9��9���9^��9���9Ό�9���99��9j��9�7�9��9x   x   �P�9
2�9�&�9�k�9���9���9� �9���9���9$�9���9���9*l�9`&�9B1�9P�9��9յ�9���9ރ�9���9��9�p�9�p�9:��9g��9��9��9L��9���9x   x   g��9�T�9G��9��9BX�9�'�9-m�9.�9�l�9�'�9�W�9��9���9-U�9���93��9LA�9;��9��9�9z�9Ch�9���9Pk�9�z�9��9-�9о�9?�9��9x   x   ���9O��9��9���9�G�9`�9X��9���9��9�H�9i��9��9��9A��9ْ�9<��9q��9���9l�9��9�v�9x3�9{/�9�u�9��9��9���9���9g��9�9x   x   �T�9h?�9��9�b�9���9��9bh�9��9a��9;a�9<��9@�9MT�9���9�;�9��9�9��9��9���9)��9"�9z��9܌�9��9��9��9 ��9�8�9%��9x   x   \n�9�9�9׀�9�j�9���9x4�93�9���9lk�9���9�9�9�m�9���9��9ؼ�9���9��9=�9��9M@�9��9��9i=�9n��9�9��9҄�9���9��9��9x   x   ~��9B��94�9�,�9Z��9���9 ��9+�9a�92��9p��9X��9U��9���9���9���9H{�9�w�9���9.�9M��9��9/��9�v�9C|�9)��9��9��9���9���9x   x   Z
�9:��9�t�9���9���9���9���9
v�9���9
�9���9���9�-�9>��9O��95��9>i�9@4�9�"�9�9��9�!�9�1�9�i�9Y��9���9��9�/�9���9���9x   x   ���9Q��9���9g��9��9�9J��9,��9���9�z�9��9���9ݝ�97�9э�9�q�9���9g0�94��9�=�9��9�1�9��9�p�9L��9l6�9J��9���9��9�|�9x   x   ���9��9�G�97W�9�X�9�G�9/�9\��9��9��9Yo�91!�9
��9݀�9��9�q�9�l�9�v�9���9��9w�9!j�9�p�9��9��9��9�"�9�q�9=�9'�9x   x   ɬ�9d�9�9슿9��9�b�9��9��9�o�9��9`j�9�-�9���9���9k��9���9|�9��9���9��9�|�9���9p��9��9���9s,�9h�9���9�o�9ι�9x   x   ��9��9�#�90#�9z�9F�9���9��92�9���9FR�9�-�9���9	7�9���9���9�9��9��9u�9���9:��9�6�9��9h,�9�T�9���92�9�9���9x   x   ���9=�9�˺9�;�9��9��9���9��9���9}��9�g�9#�95��9���9���9���9i�9���9��9n��9���9$��9i��9�"�9�g�9v��9���9��9���98�9x   x   ��9A�9��91�9|��9�e�9���9��9��9_��95q�9���9�1�9&��9��9r��9��9��9��9��9a��90�9���9�q�9���9�9��9���9*d�9q��9x   x   ���9�~�9
��9�H�9�x�9d�9v��9��9wp�9��9���9L��9��9a��939�9~��9@�9/��9A9�9k��9*��9���9��9�9�o�9��9{��9d�9�{�9�H�9x   x   㷶9*��9���9#J�9��9��9@��9(��9��9k{�9���9H��9���9��9=��9���9ǉ�9`��9���9K��9���9n��9�|�9��9u��9#��9��96��9�H�9ޙ�9x   x   },�9���9�"�9���9η9Ļ9�T�9�8�9�U�93c�9b*�9�m�9��9`��9�R�9���9�S�9���9`��9�o�9�)�9�b�9�U�9�7�9V�9�û9�η9،�9#�9���9x   x   Š�9���9�l�9Q�9S��9���9^�9��9X��9�@�9>��9�7�99*�98�9G�9H�9�6�9V*�9�6�9��9�A�9K��9���9��9���9R��9��9rl�9���9��9x   x   _"�9�l�9��9�g�9��9߿90.�9��9$�98�9��9��96e�9U��9~]�9z��9Vf�9�9���9A9�9-�9��9�/�9�߿9��9�g�9���9�l�9!#�9h��9x   x   �9��9�g�9�V�9¾9ז�9}��93��9��9�K�9�o�9��9���9���9̙�9���9���9p�9K�9���9���9j��9v��9R��9,W�9og�9��9Z��9;��9��9x   x   8ͷ9���9p�9���9��9%��9ZD�9���9�R�9�i�9���9���9+�96��9��9��9��9�h�9�T�9���9C�9��9Z�9<¾9��9特9`η9>��9W]�9���9x   x   �»9���9X޿9j��9��9��9	�9P.�9��9̏�9���9��9Ω�9'��9���9���9H��9r�9-�9��9���93��9���9�޿9���9��9���9��9�9
��9x   x   �S�9V�9d-�9��9�C�9��9���9�T�9���9 ��9e�9���9G�9f��9��9���9J��9�T�9���9%�9�B�9��97.�9��9�T�9��9~?�9���9:@�9� �9x   x   7�9���9��9|��9q��9.�9�T�9^�9T%�9ԏ�9Ĕ�9��9��9���9���9�%�9�\�9�T�9�,�9��9��9u��9}��9�5�9��9P9�9��9���9�9�9W�9x   x   CT�9��9�9��9AR�91�9���9<%�9^�95R�9H��9��9���9gQ�9i]�9w%�9X��9�
�9�S�9��9��9S��9{V�9�O�9n��9;"�9���9!�9���9�P�9x   x   �a�9�?�9�6�9K�9i�9T��9���9���9(R�9���9��9��9��9�R�9���9��9���9�i�9�H�9h8�9�?�9_�9���9$&�9\��9���9g��9���9�%�9ͯ�9x   x   �(�9ۆ�9���9�n�9U��9)��9(�9���9@��9��9�5�9��9���9��9��9��9���9�o�9#��9���9v*�9;��9۪�9��9�w�9y�9�u�9��9��9���9x   x   l�9�6�9q�9+��9V��9���9���9��9��9��9��9C�9C�9���9Z��9���9��9.�9�5�9�k�9���9S��9q!�9�D�9�`�9na�9OF�9j!�9O��9Ʀ�9x   x   ���9�(�9.d�9Ѱ�9��9���9�F�9��9"��9=��9
��9X�9BH�9s��9!�9��9�e�9!)�9 �93��9��9�A�9]��9�"�9�>�9�!�9���9�A�9���9���9x   x   ���9�6�9v��9��9ލ�9��9t��9��9�Q�9S�9*��9���9���90��9#��90��9�5�9��9�"�9���9A��9��9Us�9z��9
��9"t�9���9���9��9�"�9x   x   �Q�9F�9�\�9e��9��9���95�9_��9�]�97��9=�9���9x�9O��9]�92G�9�T�9Qo�9>s�9mJ�9���9��9p��9��9���9��9E��9�K�97s�9�o�9x   x   ~��9SG�9���9K��9��9ϋ�9-��9&�9&�9���9���9���9���9���9iG�9*��9v��9=I�9V��9z��9���9� �9 ��9C��9J �9���9��9��9�H�9'��9x   x   �R�9Q6�9f�9���9��9���9��9Z]�9:��9���9� �9���9�f�9?6�9
U�9���9��9��9���9�X�9�/�9�R�9>��9,T�9�.�9Y�9N��9��9���9d��9x   x   ��9*�9�9Gp�9Si�9$�9�U�9�U�9��9�j�9q�9F�9*�9��9p�9�I�9@�9q��9ì�9O)�9>��9���9=��9R��9a)�9Ǭ�9@��9e�9K�96p�9x   x   ��9�6�9��9�K�9uU�9�-�9���9.�9�T�9	J�9z��9�6�9N�9�#�91t�9��90��9��9���9�.�9��9�0�9���9/�9��9���9���9���9�s�9�#�9x   x   �o�9C��9�9�9>��9���9�	�9p	�9y��9q��9�9�93��9Vm�9���9��9�K�9w��9dY�9�)�9�.�9�V�9Cp�9�p�9T�9%/�9�)�9�X�9��9hL�9��9���9x   x   �)�9�A�9��9���9*D�9$��9UD�9z��9��9fA�9>,�9{��9���9׻�9.��9���9�0�9��9���9zp�9��9�p�9���9���9#1�9X��9���9y��9���9$��9x   x   �b�9ߚ�9���9s��9P��9���9���98��9;��9a�97��9F��9zC�9���9S�97�9�S�9���9=1�9Zq�9�p�9�0�9���9�S�9��9��9���9D�9��9���9x   x   =V�9v��9�0�9���9��9M��9�/�9]��9|X�9���9���9�#�9j��9Cu�9<��9���9���9a��9���9�T�9��9���9N��9^��9���9yu�9��9<#�9���9E��9x   x   ,8�9��9��9�¾9�þ9h�9q�9�7�9
R�9U(�9R��9�F�9�$�9���9��9���9�U�9���9#0�9�/�9;��9.T�9���9��9"��9%�9H�9Ӆ�9(�9ES�9x   x   �V�9l��9��9gX�9�94��9kV�9��9���9���9�y�9;c�9�@�91��9���9 �9)0�9�*�9��9�*�9�1�93�9���94��9#A�9�b�9kx�9r��9��9s	�9x   x   QĻ9%��9�h�9�h�9\��9�»9b�9];�9c$�9��9_{�9�c�9$�9Bv�9��9���9�Z�9��9���9tY�9���9!�9�u�9%�9c�91|�9���9�%�9.:�9��9x   x   BϷ9��9���9#�9�Ϸ9#��9TA�9��9���9���9x�9�H�97��9���99��9���9���9���9��9���9e��9��9A��9 H�9gx�9��9���9���9�C�9g��9x   x   \��9m�9�m�9��9���9K�9���9���9#�9��99��9�#�9�C�9���9�M�9���9�9��9���9M�9��9PD�9I#�9���9U��9q%�9���9���9�9���9x   x   �#�99��9�#�98��9�^�9v�9�A�9�;�9���9�'�9��9[��9���9���9�t�9OJ�9���9L�9�t�9l��9��9#��9��9�'�9���9�9�9�C�9��9_�9罳9x   x   0��9u��9��9ݽ�9��9O��9k�9��9TR�9���9���9���9���9m$�9q�9b��9k��9�p�9)$�9:��90��9���9��9�R�9	�9u�9��9P��9½�9驱9x   x   �9M.�9��9'�9Gױ9u��9\&�9N$�9�U�9�{�9�T�9Ԁ�9X��9w/�9�;�91��95>�9/�9���9���9[S�9�z�9#W�9�"�9�(�9���9�ֱ9q�9���9&.�9x   x   .�9JN�9ǂ�9^ͯ9��9�Ҹ92?�9�
�90��9��9Ž�9�J�9��9p�9A��9ɱ�9n�9w��9�J�9V��9ۆ�9���9a�9B>�9�и9�9�̯9(��9UP�9�-�9x   x   ���9���9�9���9�Ķ9��9!��9�K�95��9=��9�X�9�'�9���9M��9�W�9-��9���9&�9�X�9H��9���9nI�9���9���9�Ŷ9��9��97��9���9$m�9x   x   _�9�̯9z��9T�9�L�9�9���9���9i��9&�96��9�9�0�9�G�99G�9�0�9g�9��9��9���9���9#��96�9�L�9��9ό�9�̯9Q�9��9��9x   x   ?ֱ9�9kĶ9WL�9�D�9��9��9��9~��9N��9��9��9V��9��9[��9��9��9��9���9���9�9|��9�E�9�L�9BŶ9��9�ֱ9Z��9��9v��9x   x   '��9�Ѹ9D��9��9Ƙ�9;|�9qn�9�Q�9r��9
��9�m�9��9���9���9u�9�m�9R��9���9�O�9\n�9G~�9���9	�9$��9Ѹ9O��9Q"�9X�9OY�9�!�9x   x   �$�9�=�9#��9���9�9;n�92��9���91��9�G�9��9�8�9Ӛ�9y7�9?�9@G�9M��9���9��9�m�9��9R��95��9�=�9�%�9X��9^��9�K�9y��9-��9x   x   �"�9Y	�9cJ�9���9}��9�Q�9���9Ɋ�9��9r|�9���9�S�9�T�9ڹ�9C|�9)��9��9n��9�O�9���9��9I�9��9�!�90��9m��9/�9o�9��9U��9x   x   &T�9���9��9c��9ž�9���9���9Ϻ�9.?�9�p�9�3�9nm�9�2�9�o�9r@�9l��9f��9"��9(��9���9���9��9qU�9��9�)�9���9�n�9g��9)(�9*�9x   x   �y�9`��9۽�9�9���9���9SG�9K|�9�p�9�,�9d��9q��9�-�9�p�9�z�9-G�9���96��9��9(��9l��9Ew�9��9���9��94N�9M�9���9���9���9x   x   �R�9��9eW�9��9H��9m�9��9Ҹ�9�3�9j��9��91��9�2�9߹�9V�9�k�9,��9���9�X�9,��9%S�9;��9��9K��9�q�9xl�9�q�9���9���9���9x   x   �~�9I�9>&�9�9��9�9h8�9�S�9�m�9���9D��9*n�9DT�9{6�9��9��9i�9y$�9�H�9y�9"��9|�9fd�9���9K��9��9��9�e�9��9)��9x   x   |��9r��9���90�9���9���9���9�T�9�2�94.�9�2�9kT�9f��9n��9���9�/�9���9~��95��9���9���9��9�Y�98��9���9��9Z�9i��9d��9J��9x   x   �-�9�n�9@��9$G�9��9���9�7�9��9
p�9�p�9?��9�6�9���9��9OG�9���9�l�9%+�9���9k��9�1�9Lu�9S�9k��9a��9�S�9jv�9�3�9l��9��9x   x   T:�9��9,W�9�F�92��9��9��9�|�9�@�90{�9��9��9��9�G�9vW�9\��9N>�9���9J�9���9��9�9��9�J�9���9��9��9e��9@L�9.��9x   x   ���9߰�9���9�0�9��9�m�9�G�9��95��9
H�9�l�9c�9�0�9��9���9���9�C�9N��9���9�f�9��9�*�9 ��9���9C,�9���9Ne�9>��9a��9HE�9x   x   @=�9zm�9i��9i�9b��9���9#��9 ��9{��9���9H��9f�9� �9�m�9�>�9ED�9�H�9=@�9z��9���9��9S��9�9���9P�9>��9F��9�@�94I�9�B�9x   x   Y.�9(��9&�9V��9���9���9�9� �9|��9���9B��9�%�9���93,�9]��9��9�@�9ј�9�m�9���9��9X��9���9l��9و�9Jm�9���95A�9���9���9x   x   .��9�J�9)Y�9��9x��9Q�9m��9YQ�9���9��9�Z�9%J�9���9��9GK�9x��9��93n�9�_�9(U�9� :�h :� :�U�9}_�9,o�9���9b��9�L�9��9x   x   ���9���9���9`��9̉�9�o�9�o�9W��9���9��9$��9a��9s��9��9��9�g�9u��93��9uU�9{� :�.:�/:[� :@U�9V��9	��9^i�9���9���9���9x   x   �S�9W��9���9���9x�9��9��9��9ŭ�9���9VU�9N��9��9�3�9̋�9���9��9���9� :�.:�:�.:� :Q��9��9���9$��9g5�9!��9���9x   x   +{�9F��9jJ�9f��9��9G��9M��9:K�9J��9�y�9���9��9d��9�w�9 �9a,�9׆�9���9�h :�/:�.:i :Y��9/��9�-�9��9�v�9Ǹ�9U�9���9x   x   �W�9:�9���9��90G�9��9X��9�
�9�W�9���9���9�f�9f\�9�U�9X��9��9��9?��9L :�� :4 :���9��9E��9O��9iV�99\�9qh�9L��9��9x   x   w#�93?�9>��97N�9�N�9$��9/@�9P$�9I�9T��9��9���9���9���9�L�9���9���9��9�V�95V�9��9���9o��9�N�9M��9���92��9��9��9��9x   x   )�9�Ѹ9�ƶ9��9Ƕ9"Ӹ9>(�9���9L,�9ф�9^t�9��9���9��9���9.�9I�9���9�`�9d��9{�9p.�9���9b��9���9ض�9�t�9���9+�9;��9x   x   ��9�9b��9Z��9Z�9_��9���9霿9T��9�P�9Jo�9ζ�9���9UV�9	�9���9=��9�n�9�p�9��9]��9X�9�V�9���9��9�n�9�P�9ʛ�9u��9鏺9x   x   �ױ9�ͯ9,�9Lί9}ر9M$�9���9��9!q�9�O�9�t�9ݙ�9�\�9y�9���9�g�90��9���9��9Pj�9͋�9>w�9k\�9>��9�t�9�P�9q�9��9Y��9�"�9x   x   
�9���9Q��9��9���9Z�9�M�9��9��9)��9R��9wh�9���9%6�9���9C��9vB�9�B�9|��9s��9�5�9��9�h�9җ�9i��9���9��9�J�9�[�9~��9x   x   ��9�P�9���9�9��9[�9p��9=��9w*�9��9"��9I!�9���9���9WN�95��9�J�9��9�M�9)��9s��9i�98��9E��9�*�9"��9��9�[�9k�9��9x   x   b.�9".�9�m�9��9���9"#�9�9E��9B�9֝�9���9j��9s��9���9���9�F�9D�9���9���9	��9���9���9���9l�9���9f��9="�9��9a�9�n�9x   x   5B�9��9�/�9䫥9�i�9VB�9��9�.�9���9F>�9�Y�9���9��9�$�9_��9�t�9U��9�#�9��9���9WY�9>�9���9T-�96�9�D�9�h�9ݫ�9�,�9��9x   x   ��9�d�9-�91��9��9N�9��9E��9���93��9���9:{�9 ��9� �9��9���9���9\��9�|�9��9��9ћ�9��9 ��9��9J�9���9#�9pg�9��9x   x   _/�9��9�2�9^�9~x�9�V�9���9�G�9���9��9t��9�J�9.��9���9Q��9���9��9H�9؝�92�9���9{F�9���9�W�9z�9�^�9%1�9��9�,�9s��9x   x   ���9���9�]�9V��9Ԯ�9�X�9�U�9�j�90Q�9˾�9�}�9�I�9��9�A�9�@�9���9!K�9��9_��9�N�9vk�9"W�9�W�9���9Ĥ�9�^�9���9���9N��9 ��9x   x   `h�9� �9�w�9y��9���9�վ9W�96��97��9�9�l�9�R�9;&�9��9�&�9oS�9k�9L��9���9"��9�T�9�־9���9ݮ�9z�9o��9�f�9�ݨ9�^�9�ݨ9x   x   �@�9�9V�9X�9Zվ9���9C}�9�,�9���9�V�9JZ�9���9"��9c��9���9�Y�9�X�9ډ�9++�9�~�9��9�Ծ9X�9JU�9r�9}C�9Fp�9��9ね9�o�9x   x   ��9���9z��9�T�9�V�9}�9���9J��9��9��99K�9���9�5�9��9�K�9�9\�9:��9q��9a}�9V�9[U�9綼9��9��9F
�9�ݳ9�u�9�ڳ9��9x   x   �,�9���9"F�9si�9x��9�,�9��9��9a�9��9L�9��9]��9>�9p��9`�9w��9֑�9h+�9M��9j�9�D�9���9�-�9�^�9��9\��9���9��9�^�9x   x   >��9���9*��9P�9R��9��9��9�`�9ad�9���9w��9��9Ҿ�9���9�f�9b�9=�9���9���9wO�9j��9֚�9���9[-�9c�9g�9T*�9Oh�9��97.�9x   x   �;�9 ��9>�9���9ђ�9PV�9�9Ǚ�9���9\��9h+�9-,�9���9���9m��9��9�W�9��9
��9�9���9&<�9Z*�9�Q�9���9X��91��9��9�S�9M(�9x   x   :W�9���9М�9m|�9�k�9�Y�9�J�9+�9q��9k+�9lG�9+�9&��9��9�L�9�W�9�k�9	~�9ɝ�9���9�U�9G��9���9'f�9vM�9:?�9&O�9d�9��9;��9x   x   (��92y�9 I�9�H�9�Q�9	��9=��9��9��9O,�93+�9?�9%��9���9�9]S�9~H�9�F�9�y�9���9��9
l�9r��9&�9�)�9(*�9"�9��9�m�9��9x   x   U�9;��9���9���9�%�9Ѝ�9�5�9|��9��9ϵ�9i��9U��95�9v��9`&�9#��9���9���9<�9�G�9vx�9ߊ�9FX�9(��9��9'��9�Y�9���9�x�9�J�9x   x   �"�9���9���9
A�9���9@��9��9��9��9���9j�9��9���9d��9ZA�92��9���9�!�9�J�9"g�9�M�9���9G��9Ս�9���91��9.��9�O�9Se�9H�9x   x   ���9���9R��9@�9U&�9׀�9[L�9
��9�g�9/��9^M�9��9�&�9�A�9m��9���9���9#��9���9��9� �9�93:�9_��9T:�9,�9� �9���9���9���9x   x   *s�9���9���9d��9�S�9�Y�9��9
a�9c�9��9�X�9\T�9���9���9��9s�9,��9��9�{�9���9��9���9��9��9ڪ�9*��9���9�{�9���9���9x   x   .��9���9���9;K�9}k�9]Y�9X�9���9��9Y�9�l�9�I�9���9s��9.��9���9���9=k�9<��9���9�A :T):x:�(: A :���9?��9�k�9P��9���9x   x   #�9���9H�9R��9��9��9���9\��9f��9���9��9DH�9��9�"�9+��9ç�9�k�9���9���9��:�":��:	�:�#:D�:���9���9]l�9���9 ��9x   x   9�9�|�9;��9#��9���9�,�9��9?-�9���9��9П�9�{�9�9nL�9Q��9�|�9��9\��9#M:u+:�U:z�:�S:U+:�L:���9���9Q|�9���9PK�9x   x   ���9h��9��9�O�9��97��9L�9f��9�Q�9n�9 ��9
��9'J�94i�9���9��9ɩ�9C�:�+:��:��:P�:�:�+:�:}��9(��9a��9(g�92M�9x   x   �Y�9���9���9�l�9SV�9��9NX�9�l�9���9���9�X�9R�9{�9-P�9�"�9��9�B :�#:�U:�:�*:ɲ:�T:$:�B :���9#�9�R�9�z�9��9x   x   �>�9���9�G�9�X�9�ؾ9�־9�W�9VG�9���9?�92��9�n�9�9D��9�	�9ͪ�9G*:W�:�:��:�:��:/�:�):���9g
�9o��9���9�n�9*��9x   x   s��9)��9��9?Y�9�9WZ�9{��9_��9���9~-�9̖�9���9d[�9B��9�<�9���95y:��:�T:��:�T:U�:y:���9:�9���9%\�9���9g��9�*�9x   x   +.�9O��9kY�9˰�9
��9�W�9ǆ�9�0�9x0�9U�9xi�9��9x��9���9U��9Ǧ�9�):�$: ,:\,:g$:�):Ч�9���9���9���9�9Wg�9#W�991�9x   x   �9:�9
|�9���9F|�9��9��9�a�9��9��9�P�9�,�9b�9��9g=�9���9?B :N�:�M:��:7C :1��9�:�9ґ�9T�9Z.�9S�9���9M�9wa�9x   x   �E�9��9 `�9L`�9� �9�E�9�9�"�9Qj�9���9�B�9�-�9���9}��9>�9 ��9���9���9J��9���9���9�
�9���9���9V.�9<@�9���9 i�9^$�9]�9x   x   Qi�9���9�2�9L��9i�9�r�9:�9G��9�-�9z��9�R�9��9?]�9f��9�#�9���9���9���9z��9^��9�#�9���9h\�9�9�R�9���9�.�9냺9�޳9rq�9x   x   ���9%�9.�9��9uߨ9́�9^x�9P��9Zk�94��9[g�96��9Ԋ�9S�9ʿ�96~�9�m�9%n�9�}�9g��9pS�9���9���9Fg�9���9�h�9Ӄ�9Tw�9U��9��9x   x   \-�9>h�9.�9Ą�9Q`�9�9Zݳ9z"�9��9�V�9��9�p�9�{�9!h�9O��9ʦ�9<��9>��9���9�g�9({�9�n�9<��9�V�9��9�#�9m޳9(��94]�9���9x   x   ��9i�9V��9V��9&ߨ9�q�9�92a�9�0�9
+�9���9@�9dM�9�J�96��9x��9L��9M��9 L�9�M�9��9���9I*�9�0�9�`�9��9�p�9!�9m��9y��9x   x   �	�9,�9�p�9v��9�i�9�b�9tq�9i?�9ei�9��9�2�9�9И�9���9���9��9���9N��9x��9 �9�3�9���9$j�95>�9�q�9�e�9g�9�9Qo�9���9x   x   ���9sx�9��9�q�9,��9桫9ؚ�9&�9���9�.�9���9"��93.�9;��9I��9���9���9f0�9 ��9��9�-�9���9?�9���9՞�9���9�s�9Ͻ�9y�9��9x   x   p�9���9ck�9�|�9	��9���9�z�9G��9���9��9��9���9���9V��9���92��9���9���9H��9&�9��9)��9�x�9U��9௨9G}�9�g�9&��9�p�9���9x   x   X��9�p�9{|�9���9֭9H��9���9.\�9��9W7�9��9
��9��9���9o��9e��9��9G��9<8�9���9pZ�9���9���9g֭9M��9�}�9u�9���9�<�9s=�9x   x   4h�9��9J��9�խ9/ų9�'�9a��9�{�9B��9�y�9�;�9k��9B�9~��9��9���9:�9�x�9��9�|�9���9�(�9�ĳ9�խ9(��9y}�9�e�9�}�9bҞ9�{�9x   x   !a�9`��9���9���98'�9k��9��9,��9��9B��9j��9�9+s�9�t�9��9i��9��9o�90��9���9V��9�&�9���9Ѿ�9Ҡ�9.d�9'�9g	�9�
�9�&�9x   x   ;o�9 ��9Hy�9w��9���9���9��9���9L�9h��9��9�u�9��9�r�9	��9]��9�H�9���9q�9���9���9���96y�9ݗ�9�n�9��9٬�95�9���9��9x   x   �<�9�9���9�Z�9�z�9���9���9���97/�9���9���9.��9��9%��91��9{/�9���9i��9ۺ�9/y�9�Z�9q��9��9�=�9��9���9���9#��9��9��9x   x   �f�9���9���9n��9:��9@�9�K�9/�9��9��9���9�9���93��9ۚ�9s0�9H�9T�9���9k��9���9���9�d�9���9�*�9<Q�9��9�S�9�)�9��9x   x   ��9E,�9��9�5�9�x�9���9��9m��9��9��95<�9�<�9ͣ�9d��9���9���9���9v�9q7�9�9�,�9���9i:�9�<�9^��9�7�9�4�9"��9>�9�9�9x   x   �/�9��9��9���9�:�9���9��9���9}��9;<�9$z�9�;�9 ��9���9��9���9�:�9C��9r��9���9�-�9���9�P�9��9C��9���9q��9�
�9 P�9a��9x   x   �9���9��9���9w��9��9Cu�9.��9&�9�<�9<�9��9���9�s�9��9;��9���9S��9��9��9�s�9��9�U�9W��9���9o��9��9�W�9���9�q�9x   x   ��9�+�9"��9���9r�9�r�9��9F��9��91��9s��9���9��9Tt�9<�9���9k��9�,�9=��9��9`��9#��9d��9���9���9���9��9A��9���9��9x   x   ��9+��9Ԏ�9���9���9�t�9"s�9���9Ƀ�9��91��9�s�9�t�9���9���9��9j��9̊�9�:�9���9/(�9!�9��9[;�9�;�9��9-!�9)�9���9~8�9x   x   ��9���9e��9Ă�9x�9��9���9���9���9���9��9��9��9��9��9���9���9K��9�O�9���9+��95A�9���9C�9<��9G@�9��9���9�R�9,��9x   x   ��9P��9n��9��9���9	��9E��9�0�9�1�9��9ف�9]��9���9���9L��9���9���9n��9��9���9%:�\:�:�:�]:�$:���9f��9O��9޵�9x   x   ���9���9W��98��9�:�9��9J�9g��9�I�9���9m<�9���9���9���9y��9+��9���97��9�?:h�:oj:|�:��:h�:�j:��:�?:��9B��9��9x   x   a��9�/�9Ü�9���9�y�9��98��9O��9Y�93x�9P��9X��9�.�9l��9���9Y��9���9��:r�:�N:�	:�	:��	:�	:7O:��:�:M��9���9���9x   x   ���9 ��9���9%9�9q��9��9u�9��90��9�9�9���9���9���9�<�9VQ�9t��9E@:��:�:�K
:P�:jE:j�:�J
:s�:`�:�?:
��9�T�9=�9x   x   �9���9�9��9@~�9���9��9�{�98��9�9���9v�9� �9M��9(��9���9$�:O:�K
:�`:v{:{:Jb:hL
:kN:�:%��9���9	��9�"�9x   x   44�9�.�9L��9\�9���9���9O��9�]�9��9�/�9:1�9�v�9���9*+�9���9N&:hk:�	:��:�{:�:{:��:m	:�k:�%:���9V.�9��9�u�9x   x   ���9���9���9���9#+�9Z)�9���9���9,��97��9���9���9���9j$�9WD�9O^:��:��	:F:y{:�{:aG:��	:{�:_:mE�9L"�9-��9F��9Ĭ�9x   x   k�9��9�z�9���9.ǳ9m��9Z|�9R�9h�9.>�9�T�9�Y�9=��9{��9	��9q:�:��	:J�:�b:��:�	:��:�:���9ń�9���9[�9�U�9�<�9x   x   H?�9N��9'ï9�ح9Uح9���9%��9}A�9x��9�@�9��9v��9���9K?�9�F�9�:�:#	:�K
:(M
:�	:ǌ::;G�9&@�9`��9b��9��9�A�9{��9x   x   s�9N��9���9���9Ʊ�9ϣ�9,r�9��9�.�9r��9{��9���9���9�?�9��9�_:9l:�P:��:<O:Fl:m_:���9N@�9G��9��9��9x��9�-�9��9x   x   �f�9��9#�9��9��9 g�9U�90��9U�9�;�9$��9���9ދ�9��9#D�9g&:=�:�:t�:��:&:*F�9+��9���9��9���9,;�91U�99Q�9x   x   h�9u�9�i�9'w�9Xh�9�)�9��9=Ĵ9��9�8�9���9J��9&��9.%�9���9���9A:P�:�@:���9���9�"�9���9x��9���9;�9��9�ô9��9*�9x   x   ���9���9���9���9��9�9�8�9�ô9kW�9���9��9�[�9/��9�,�9q��9���9���9���9ƈ�9���9+/�9���95[�9��9A��9�T�9�ô9�9�9��9��9x   x   �o�9z�9Hr�9B>�9�Ԟ9F�9���9 ��9Z-�9�A�9�S�9���9S��9W��9�U�9��9���9p��9 V�9���9���9c��9zU�9A�9r-�9x��9���9��9WӞ9?�9x   x   G�9���9���9�>�9�}�9�(�9i�9v�90��92=�9ǭ�9Pu�9� �9�;�9��96��9ն�9��9	>�9H#�9�u�9���9&<�9ǋ�9�9��9])�9o�9�>�9粖9x   x   6�9uE�9�\�9�f�9�C�9���97r�9�9f(�9�K�9���9�r�9;y�9y��9�W�9���9[�9��9�w�9�o�9���9N�9+)�9��9�q�9���9@�9�e�9]�9aE�9x   x   E�9FH�9m�9�Ò9�9뢢9�J�9�9��9R�9o��9� �9���9�l�9���9���9�m�9a��95"�9���9�P�9w�9���9XL�9���9��9eƒ9h�9�F�9�B�9x   x   �[�9�9��9���9�9���9��9�ĺ9�v�9ܻ�9q�9	�9IS�9���9?��9"��9�Q�9��9R�9ҹ�9�w�97Ǻ9�9ᱧ9��9۬�9��9��9[`�9_s�9x   x   ee�9Ò9?��9|�9�Z�9ѣ�9���9p��9L�9�p�9���9n$�9�(�9�*�9�,�9'�9�%�90��9Kr�9N�9��9̀�9��9�[�9��9���9�ǒ9c�9뷍9f��9x   x   �A�9��9&�9#Z�9�~�9Y�9��9a��9�^�9�K�9�'�9���9H�9�0�9F�9��9$&�9�J�9[\�9���9ԃ�98Z�9k}�9�Y�9��9G��9�@�9���9�+�96�9x   x   E��9��9H��9�9�X�9���9���9���9�~�9h3�94��9��9f��9���9��9��9_6�9_��9���9���9���9Y�9���9⯧9ܢ�9���9F�9���9���9g�9x   x   �o�9�H�9� �9��9V��9P��9��9r�9/{�9N��9|v�9Ɵ�9�c�9j��9�v�9c �9�v�9`�9�	�9T��9���9�}�9	�9lG�9o�9ə�9�ۣ9�C�9hݣ9"��9x   x   �9e��9�º9���9V��9��9,�9���9�)�9ӊ�9���9.�9/�9r��9���9+�9��9��9r��9��9B��9ĺ9���9=�9�Q�9z�9���9���9�w�9hR�9x   x   %�9�9Pt�9IJ�9�]�9~�9�z�9�)�9<�9.��9��9+��9l�9���9�:�9�*�9x�9�97\�9�J�9�u�99�9�$�9ջ9% �9D"�9θ9�$�9�!�9�ӻ9x   x   eH�9+O�9y��9�n�9FJ�9~2�9���9���9��9��9=��9`��9"�9���9e��9S��9�4�9wH�9r�91��9,O�9�K�9��9�h�9���95�9$3�9ە�9�h�9���9x   x   ��9j��9	�9���9�&�9T��9v�9���9��9N��9��9��9��9��9�w�9k��9�%�9p��9�9���9���9^+�9���9oj�9�<�9�2�9*?�9�j�9@��9�,�9x   x   o�9��9��9�"�9׊�9�9~��9x.�9_��9���9;��9���9/.�9_��9b�9܋�9�$�9d�9��9mm�9���9Xj�9���9�^�9ٗ�9b��9]]�9B��9�h�9���9x   x   �u�9��9$Q�9'�9G�9���9�c�9Z/�9��9��95�9s.�9le�9���9�G�9�#�9�O�9���9ss�9�C�9��9t��9���9��9�9���9���9.��9(�9�@�9x   x   \��9dj�9؝�9�)�9o0�9���9���9��9b��9Y��9���9���9��9].�9�+�9,��9�i�9��9���9��9_��96j�9i-�9Y�9��9!.�9�i�9u��9#�9���9x   x   U�9���9Ը�9,�9�E�9�9bw�9|��9�;�9���9�x�9_�9YH�97,�9o��93��9U�9%�9���9�9�9Ĉ :$:��:RD:�:D:Ɖ :�5�9���9��9x   x   C��9#��9;��9�&�96��9���9��9q,�9�,�9� �9���9K��9%�9��9���9���9���9��9�:c/:a:`�:�:��:��:�_:�0:V�:@�9���9x   x   UY�9�l�9wQ�9<&�9�&�9�7�9Bx�9���9z�97�9�'�9�&�9�Q�9fk�9#V�9`��91j�9	 :z:/q	:׹:�(: �:i':K�:Bp	:ly:U :`k�9g��9x   x   ۊ�9���9�9��9�K�9��9k�9�9���9K�9���9��9��9ۍ�9��9	�9O :�<:_:�:�B:ad:�e:B:N:�:�<:� :S�9"�9x   x   w�9G"�9��9s�9^�9���9
�9@��9#_�9u�9�9�"�9>v�9~��9���9�:�z:�:�:(�:�:^:\�:F�:��:#:z:��:��9p��9x   x   �o�9
��9���9�O�9"��9��9C��9;��9�M�9���9Y��9�p�9�F�9��9U<�9�0:r	:h:z�:3�:K�: �:��:9�:�:Zr	:m1:;�9i�9OG�9x   x   ���9�Q�9\y�9��9W��9���9ʆ�9͇�9�y�9S�9��9���9��9��9r� :�b:�:�C:��:��:~�:]�:��:}D:x�:�a:1� :���9��9���9x   x   �N�9��9ɺ9��9 ]�9�\�9>��9�Ǻ9Y�9�O�9�/�9�n�9̯�9in�9:�:8*:�e:�^:��:��:M`:=f:�(:��:�:l�9���9�n�9�.�9x   x   ?*�9I��9�9���9o��9i��9��9���9")�9z��9L��9���9���9 2�9��:��:ԧ:�f:v�:m�:-�:tf:ʧ:߽:��:�2�9 �9���9Ӳ�9>��9x   x   ��9N�9��9�^�9�\�9w��9WK�9��9�ٻ9�m�9po�9d�9(��9;�9�F:�:J):�C:��:.�:%E:_):�:gF:��9���9�c�9n�9�m�9Nٻ9x   x   s�9q��9��9��9��9���9s�9V�9�$�9���9�A�9��9�$�9��9c�:��:=�:�:�:�:3�:��:��:�9�%�9U��9�C�9��9�$�9'W�9x   x   ��9G�9��9?��9[�9B��9���9a~�9�&�9:�9)8�9���9 ��9=3�9�:�a:7r	:z	:u	:cs	:eb:h:o3�9"��9j��9�5�9�9�9\(�9�}�9���9x   x   AA�9
Ȓ9/��9ʒ9�C�9��9}ߣ9M��9�Ҹ98�9:D�9�b�9���9�n�9� :3:F{:>:R{:]2:֊ :�l�9i �9�c�9�C�9�9�9)Ҹ9=��9�9
�9x   x   �f�9� �9c�9ke�9���9ˮ�9�G�9���96)�9���9ho�94��9��9(��9:�9L�:	::Æ:�<�9���9��9���9�m�9қ�9(�9��9!I�9���9���9x   x   �]�9H�9�a�9���9$.�9���9��9^{�9�%�9Mm�9ͯ�9$m�9��9o�9���9��9Qn�9�	�9���9��90�9�n�9���9�m�9 $�9k}�9�ߣ9e��9.�9R��9x   x   �E�9�C�9�t�9#��9l��9�92��9�U�9`׻9���9�0�9���9�D�9G��9��9���9���9��9���9�G�9���9�.�9���9vػ92V�9���9?	�9=��9��9�u�9x   x   �3k9��m9��t9S��9/��9@Β9)v�9�P�9�˸9sH�9�7�9c��9���98�9k��9�h�9���9�4�9���9k��9�7�9!K�9͸9�P�9�t�9�Β9���9끀9a�t9�m9x   x   �m9�[r9r�{9І�93>�9���9�+�9{��9�d�9w��9#u�9"��9ڷ�9k�9#_�9�[�9[m�9��9r��9�w�9���9�b�9��9�,�9��9�?�9|��9h�{9�Zr9�m9x   x   ��t9m�{9!�9Dk�95d�9Ѻ�9m�92Ҵ9���9=��90
�9��9.�9h�9v�9b�9�9���9��9���9I��9�Դ9T�9r��9b�9Ak�9��9t�{9<�t9~�r9x   x   ���9���9�j�9��9O�9J�9Y��9���9e�9�J�9b��9���9���9NF�9QI�9���9���9� �9_K�9�f�9&��9|��9T�9s��9}��9$k�9���9�~�9{�|9��|9x   x   ��9�<�9 c�9��9B��9�(�9��9=�9�q�9g�9�(�9���9���9��9���9���9Q&�9&�9%p�9a�9d�9a)�9)��9:�9�b�9�:�9���9+�9���9L�9x   x   �˒9���9;��9H�9n(�9m�9Ծ9��9��9J��9e�9�[�9�d�9-e�9�\�9%d�9Z��9���9;��9?Ծ9o�9�*�9Z�9���9?��9�˒9���9�ݍ9�ݍ9�9x   x   �r�92)�9e�9鸯9��9�Ӿ9e��9��9ƶ�9�V�9���9�F�9`/�9�F�98��9X�9���9�9��9?Ծ9�9���9��9�(�9Or�9��9s�9y,�9��9b�9x   x   �L�9|��9�ϴ9���9��97��9j�9w��9�J�9ߛ�9?��9] �9��9"��9'��9,K�9���9}�9щ�9��9 ��9Ѵ9���9�L�9_��9���9F��9��9۷�9j��9x   x   ȸ9Na�9ѥ�9�b�9Sp�9"��9D��9�J�9OG�9�C�95�9��9��9�C�9F�9�K�9���9Щ�9�m�9c�9o��9_�9�ȸ9a�9�ֳ9���9#�9���9�׳9U�9x   x   3D�9���9\��9PH�9� �9S��9`V�9���9�C�9�%�9^ �9N!�9@%�9�D�9���9V�9���9� �9�K�9P��9��9�F�9@�9���9ڴ�9Z3�9P2�9��9��9�B�9x   x   �3�9yq�9B�9(��95'�9d�9+��9��9C�9m �9Ce�9f �9��9ώ�9���9�b�9M%�9���9F�9^t�9�2�9;N�9���9�S�9%�90�9�'�9�T�9���9�O�9x   x   ��9���9O��9���9c��9�Z�9UF�9c �9X��9�!�9� �9���9��9�D�9�[�9��9U��9o��9/��9���9�h�9!�9۽�9F�9���9���9�C�9��9�9�g�9x   x   ���9t��9��9��9���97d�9q/�9@ �9]�9�%�9�9��9�1�9�c�9���9U��9��9ε�9���9U��9�*�9�2�9H��9O��9�3�9>��9��9�2�9Q,�9���9x   x   I4�9h�9?�9�D�9T�9e�9	G�9��9�D�9�E�9���9�E�9Vd�9z�9G�9��9�g�9�3�92�9v/�9���9l��9t� :$:#:�� :$��9/��9�1�9y1�9x   x   ��9�\�9lt�9yH�9}��9-]�9+��9l��9�G�9|��9g��9]�9���9�G�9�p�9o[�9o��9���9�E :Q
:`n:�K:�:��:܀:�K:zo:	:>F :��9x   x   �e�9�Y�9R�9Z��9"��9.e�9�Y�9�L�9�M�9%X�9�d�9���9���9��9\�9�f�9�9*�:W�:T�	:��:��:��:�:��:�:8 
:x�:"�:��9x   x   ���9l�9��9 ��9R'�9��9���9'�9��9��9�'�9���9��9�i�9���9��9=�:|:��:��:�}:�R:�:BQ:�:]�:��:�{:�:��9x   x   3�9F��9͗�9��9��9٬�9��9]�9��9��9���9i��9���96�9r��9��:}|:5�:d�:�v:�7:ާ:-�:j7:&v:m�:v�:�|:��:��9x   x   ���9���9y	�9�L�9Mr�9��9%��99��9�q�9>O�9��9՚�9��9<5�9BG :m�:��:ɖ:�y:�;:��:+f:��:;:�z:��:��:F�:�G :8�9x   x   a��9�x�9��9�h�9��9a׾9�׾9��9;g�9���9�x�9%��9v��9M3�9
:� 
:ԛ:_w:�;:��:6\ :d[ :;�:�;:|v:�:?
:�:0�9r��9x   x   l8�9��9.��9���9r�9�9��9Z��9��9���9�7�9~m�9�/�9!��9vp:m�:�:�8:��:�\ :�R!:i\ :M�:}9:�:��::p:O��9q1�9�l�9x   x   "L�9`d�9�ִ9X��9�,�9s.�9ܺ�9�մ9	d�9�K�9�S�9��98�9���9N:��:�T:`�:Og:\ :�\ :�g:)�:�S:��:'O:��9F5�9o �9$S�9x   x   vθ9"��9��9t�9ӣ�9|�9��9���9�͸9 F�9o��9���9��9K� :ǃ:e�:.�:��:�:@�:�:n�:��:��:�:{� :���9Z��9���9�E�9x   x   R�9�.�9&��9���9��9�9Z-�9�Q�9��9��9�Y�9VL�9���9':��:��:�S:g9:�<:/=:P::dT:��:T�:': ��9�K�9�Y�9���9E�9x   x   �v�9@��9�d�9���9�f�9���9!w�9���9:ܳ9��9b+�9��9l:�95&:ރ:y�:#�:<x:Q|:�w:��:;�:f�:/':�<�9V��9�,�9N��9�۳9���9x   x   �В9�A�9�m�9]n�9n>�9В9��9���9K��9p9�9��9&��9���9Ô :�N:��:Ҝ:��:`�:̝:��:�O:͔ :`��9g��9`�9�8�9*��9��9��9x   x   /��9y��9H"�9͊�97��9߉�9 �9p��9�(�9I8�9�-�9*J�9v��9H��9dr:�
:��:s�:�:o
:q:��9;��9L�9�,�9�8�9�(�9���9��9>��9x   x   !��9ш{9�{9���9���9��9�0�9	��9癲9̸�9�Z�90��9�8�9���9�:�:~:�~:��:�:���9�5�9���9}Y�9���9Й�9���9+2�9�9:�9x   x   �t95]r9��t9e�|9���9}�9��9x��9�ܳ9<��9��9��9�1�9�6�9�H :M�:��:*�:�H :v1�9>2�9� �9;��9��9۳9Y��9V�9���9���9o�|9x   x   ݢm9��m9��r9�|9��9��9�9���9��9�G�9�T�9�l�9���96�9��9x�9��9S��9�9�90��9�l�9�R�9.E�9A�9`��9��9E��9x��9��|9W�r9x   x   x�B9��E99�N9|�\9�Hp9l9�9C�92��9���9@U�9�9�^�9'c�9���9�N�9�9�9EO�9]��9�c�9^�9��9�W�9F��9��9�A�9�8�9XJp9B�\9NN9��E9x   x   ��E9�AK9�[V9�yf9c:{9V�9w �9=�9q�9��93��9��9��9��9���9��9��9��9�9���95��9o�9;�9��9<�9�;{9�vf9�ZV9kDK9��E9x   x   �~N9eZV9,c9Ìt9�	�9o�9��9e�9~��9�t�9��9�M�9\5�9j�9a��9��9N4�9�L�9��9�t�9P��9�f�9J�9�m�9��9�t9�c9�YV9|N9y�K9x   x   ��\9wf9v�t9�f�9�/�9vU�9�[�9?��9���9��9�b�9���9���9���9���97��9���9d�9���9���9x��9\[�9!W�9�0�9�f�9�t9�tf9��\9��W9#�W9x   x   �Cp9�6{9l�9�.�9Ș9�U�9"k�9i��9��9r��9AA�9���9x�9(��9�9���9�>�9��9� �9��9�l�9+U�9�Ř9�.�9A	�9�6{9�Ep9Œi9�Jg9m�i9x   x   >6�9��96m�9BT�9U�9s��9���9e��9��9�S�9_R�9`<�9R��9~��9�<�9�R�9�T�9���9w��9I��9	��9�V�9�U�9l�9��9]6�9�=�9�z|9P||9�>�9x   x   I?�9O��9!�9�Y�9	j�9_��9|��9֫�9.�9<�9UM�9���9q��9,��9�K�9��9��9��9��96��9�j�9MX�9h�9���9�>�9&��9Gh�9c��9Df�9���9x   x   ߪ�9��95b�9��9�9���9��9�:�9m��9�(�9Z��9��96��9h��9�(�9���9}<�9N��9.��9e��9���9�b�9/�9���9U��9���9R`�9�a�9���9��9x   x   ��9m�9H��9<��9��9ҙ�9��9?��9���9/��9��9B��9c�9���9���9_��9�9��9��9��9���9ql�9��9@[�9�Ϋ9�<�9i��9�;�9�Ϋ9-[�9x   x   %P�9���9!q�9~��9���9�R�9��9�(�9 ��9��9;f�9�g�9��9١�9�(�9��9`T�9���9���9�o�9i��9�Q�9���9`ս9���9���9���9���9�ս9���9x   x   ��9ϳ�9
��9�_�9|?�9OQ�9�L�95��9��9[f�9���9uf�9
�9'��9�L�9�P�9�=�9r_�9���9ڵ�9`�9]��9�!�9u��9�m�9�_�9�n�9��9��9=��9x   x   MY�9t�9AJ�9���9��9�;�9w��9D��9���9h�9�f�9Q��9b��9���9!<�9��9���9#J�9N�9qX�9o��94��9��9;2�9��93��9�0�9��9���9���9x   x   ^�9��9Z2�9���9O�9ݿ�9���9���9�9l�9�
�9���9���9K��9��9��9b0�9v	�9�^�9��9���9�G�9dY�9��9m%�9z��9�X�9rG�9���9p�9x   x   ��9�9��9��9���9���9Ѡ�9v��9���9.��9V��9x��9ۿ�9D��92��9 �9 �9l��9�m�9�]�9%�:��:Y:,:�:IY:.�:��:�^�92n�9x   x   �J�9���9o��9���9�9�=�9�L�9.*�9|��9�*�9WN�9�=�9��9���9��9��9�J�9�8:��:�U:�d:��:"B:��:�B:j�:@e:
V:��:8:x   x   /6�9���9��9���9M��9T�9g�9*��9���9Z�9S�9@��9���9v�9���9�6�9H:H:�:�:��:n:=d:�d:u:�:/:�:�:,H:x   x   �L�9I�9�3�9O��9?@�9�V�9N�9o?�9'�9�W�9�@�9���9�2�9�9GL�9vH:5	:�:��:�`:�:�c:�0 :Xb:�:9a:�:':H4	:�H:x   x   ���9�9NM�9Ce�9 ��9���9G��9ڮ�9՝�9���9Ic�9�M�9��9g��9�9:":b:B�:5�:d� :�Y$:�'&:F)&:ZZ$:�� :��:��:�:�:�9:x   x   c�9B�9+��9���9L#�9ʬ�9׊�9Y��97!�9m��9H��9��9�b�9�q�91�:n�:��:��:�":�&:��):e�*:��):m�&:�":��:X�:k�:��:�s�9x   x   ^�9���9|v�9D��9Q��92��9���9(��9��9)u�9��9�]�9�9{b�9�W:�:�a:c� :��&:1+:�o-:wp-: 2+:��&:�� :�b:r:*X:�a�90�9x   x   V�9�9���9���9sp�9l�9�o�9ꮴ9.��9;��9S�9t��9���9��:Eg:��:�:[$:��):dp-:ˡ.:Xp-:Q�):8[$::��:g:��:���9��9x   x   �X�9q�9Ei�9�^�9JY�9X[�9�]�9kh�9�r�9X�9���9���9HN�9/�:��:':Af:�)&:��*:fq-:�p-:a�*:�*&:$f:p:��:P�:�L�9"��9���9x   x   ���9��9g�9�Z�9@ʘ9�Z�9��9=�9-��9�ǿ9�(�9N��9�`�9]:�E:Tg:�3 :�+&:��):G3+:�):�*&:_2 :4h:sE:]:�b�9��9	(�9�ƿ9x   x   ���9[�9@q�9�4�9y3�9<q�9��9A��9�a�9�ܽ9��9�9�9Ų�9�:(�:h:We:�\$:z�&:4�&:I\$:�f:rh:��:w:���9�9�9o��9=޽9�a�9x   x   �C�9�
�9!�9�j�9��9�	�9�D�9���9�ի9���9Zu�9��9j-�9�:�F:�:�:u� :�":� :A:3:�E:�:�/�9��9[v�9���9ի9���9x   x   �:�9A{9��t9��t9�?{9�;�9��9�ƚ9�C�9A�9lg�9-��9���9=]:1�:��:Sd:^�:(�:Wd:��:X�:s]:��9)��9�g�9��95C�9�ǚ9/�9x   x   �Mp9E{f9�#c9�{f9#Np9tB�9�m�9�f�9)��9�9#v�9p8�9�`�9
�:�h:�:
�:R�:\�:�:#h:��:�c�9�9�9Hv�9��9���9�f�9�k�9�B�9x   x   �\9�^V9J_V9�\9��i9C�|9���9�g�95B�9u��9I��9���9�N�9:�:uY:�:�:�:*�:kY:��:�M�9R��9G��9K��9�B�9�f�9���9�|9=�i9x   x   c�N9�GK9��N9c�W9Rg9΄|9(k�9mǚ9�ԫ9mܽ9�&�9���9���9[e�9��:T:�6	:t:�:ac�9���9Y��9�'�9�ݽ9Eԫ9ǚ9�j�9F�|9TOg9?�W9x   x   ��E9	�E9 �K9��W9��i9eB�90 �9���9�`�9eǿ9_��9���9w�9�s�9�::dJ:zJ:%;:�u�9&�9I��9q��9�ſ9j`�95��9��9�A�9n�i99�W9t�K9x   x   �G98�92 9	�09P�G9X�d9��9b��9JG�9-�9>S�9��9�|�9���9�_:"�:_:��9~�9}��9�R�9�.�9�F�9���9I�9��d9�G9|�09� 9�9x   x   ��9_9J`)9�z<9�-U9�r9Z)�9I6�9��9�B�9�r�9e��9��9�E�9��9���9ZF�9���9��9�q�9B�9,�9f7�9|*�9$�r9-+U9Jv<9�])9�b9��9x   x   [ 9�^)9�89�wM97)g9���9 �9�*�9���9�*�9�I�9^��9f��9޸�9���9���9���9���9�K�9,�9���9+�9��9��9�,g9�xM9��89�_)91 9��9x   x   ��09�w<96vM9'Ec9XO}9�L�9"�9U2�9?��9���9��9�9�_�9%�9�$�9+`�9��9̮�9���9���93�9��9�O�9�M}9�Bc9�sM9�r<9��09|+9�+9x   x   p�G92)U9>&g9�M}9�m�9�s�985�9�9N�9���9��9-��9A��9�z�9[��9Ͽ�9̛�9>��9M�9&�9>5�9�r�9(m�9lO}90)g9U,U9�G9��?9�F=9��?9x   x   �d9��r9���9{K�9Qs�9��9��9��9�W�9��9w��9���9���9@��9*��9��9��9uV�9��9��9G��9\s�98L�9O�9�r9g�d9e[9(0V9%/V9f[9x   x   -�9�%�9O�9�9�3�9�9ƿ9�%�9�b�9g�9��9m��9�2�9���9-��9�9�c�9�$�9�ƿ9g�94�9��9.�9o'�9��9��{9ǃu9Ps9K�u9`�{9x   x   C��92�9�'�9�/�9[�9��9,%�9Ċ�98��9���9�D�9��9M��9�D�9���9���9m��9p%�9#�9`�9�/�9x'�9m1�9���9���9��9_�9!`�9��9k��9x   x   �A�9�9݄�9Z��9Y�9}V�9�a�9
��96�9?�9��9�9�9��98�9`��9�a�9V�9d�98��9���9��9�A�9�Ϥ9���9벟9��9+��9��9�Ϥ9x   x   �&�9�=�9�&�9���9���9?�9��9g��9:�9]9�9B��9���9\8�9_	�9���9�9L�9���9���9q&�9=�9'�9�ڹ9��9��9�'�9p)�95�9��9)ڹ9x   x   �L�9@m�9�E�9��9��9R��9���9�D�9��9q��9���9���9��9D�9M��9���9��9W��9=G�9�m�9�L�92��9���9*�9���9	��9*��9�)�9���9���9x   x   ���9*��9]��9;�9p��9���9D��9P��9��9��9���9��9Ͳ�9/��9M��9߽�9��9���9���9ܱ�9�^�9�H�9~R�9%�9��9���9F&�9nR�9.I�9�]�9x   x   nv�9"��9¤�98]�9��9���9�2�9��9#�9a9�9Z�9L��9�2�9z��9���9/]�9���95��9�x�9t��9��9)7�9���9�~�9��9q~�9���9G7�9Y�9���9x   x   ��9fA�9��9W#�9@z�9���9���9)F�9f�9�9�E�9L��9"��9
z�9�"�9d��9�A�9v��9�� :�:��:�E	:�:�:1::{F	:��:�:�� :x   x   .]:@��9���9�#�9v��9)��9ܠ�9֋�9a:�9��9w��9��99��9�#�9���9m��93]:H�:�T
:��:�:ɒ:a�:L*:��:�:�:D�:�S
:��:x   x   �:ު�98��9
`�9���9���9��9���9��9!�9���9���9k_�9���9N��9̒:�U:)X:�D:Σ:�:�[!:�#:�#:6\!: :N�:E:�Y:�U:x   x   z]:�D�9#��9O�9���9!�9-g�9��9�e�9<�9ܝ�9��9��9"D�9%^:}V:G�:#:�:�.$:f�(:	�+:��,:+�+:�(:;0$:#:M":��:�V:x   x   Һ�9���9m��9v��9���9�Y�9�(�9�)�9�Z�9���9���9��9W��9��9��:=Y:�#:n�:�R':��-:N'2:ۂ4:�4:g(2:"�-:WR':�:�#:�Y:��:x   x   }�9;��9M�9z��9��9� �9�˿9N �9��9-��9�L�9��9~�9� :�V
:�F::RS':G/:�g5::L9:��::\J9:�h5:"H/:�R':&:�F:V
:&� :x   x   |��9�r�9\.�9 �9C�9���9���9-��9Y �9�,�9dt�9A��9���9�:Q�:�:�0$:�-:Lh5:V�::�=:p�=:1�:::g5:c�-:�0$:¥:�:��:ζ�9x   x   �S�9D�9���9�6�9�9�9���9�9�9A6�9Ƌ�9D�9�S�9f�9�9?�:E�:�":��(:4)2:M9:��=:�S?:��=:;N9:�(2:��(:�":�:��:�9�f�9x   x   �0�9��9�.�9G�9�w�9'y�9:�9[.�9�9�.�9:��9)Q�9X?�9�I	:��:7_!:�+:R�4:֤::��=:R�=:��::�4:��+:�^!:��:J	:�@�9�P�9u��9x   x   �H�9_:�9v�98T�9�r�9LR�9��9�8�9`I�9��9Y��9d[�9���9*:��:�#:S�,:چ4:�L9:��::EO9:Y�4:y�,:�#:�:::B��9K[�9���9h�9x   x   ���9�-�9��9RW}9rZ}9���9N.�9#��9�פ9M��9F3�9�.�9:��9Z:�.:�#:��+:�+2:Xk5:<i5:1*2:M�+:#:�.:�:��9B/�9!2�9ƈ�9�ؤ9x   x   ��9��r9�4g9.Lc964g9��r9��9l��9���9���9o��9���9��9 :y�:�`!:�(:��-:�J/:��-:9�(:�_!:h�:&:��9���9���9���9���9���9x   x   `�d9b1U9��M9}M97U9��d9�{9$�9C��9�0�9���9|��9}��9�:��:�$:34$:�U':NU':3$:v$:��:�:_��9���9���9�1�9��9$�99�{9x   x   d�G9�{<9�89�{<9J�G91([9�u9�f�9�9D2�9��9�/�9T��9HK	:��:��:�!:=�:�!:��:b�:�J	:��9x/�9���9�1�9��9�g�9��u9�&[9x   x   ��09�b)9�e)9��09_�?9�:V9�\s94g�9���9���9�2�9�[�9�@�9��:��:�H:�%:�&:�H:��:��:�A�9�[�9�1�9W��9���9ag�9}\s9N<V9�?9x   x   ! 9�f9s 9D+9<O=99V9֍u9	$�9f��9���9��9�Q�9��9��:~W
:�\:��:\:�W
:��:H�9
Q�96��9�9���9�"�9 �u9d;V9eQ=9�+9x   x   D�9\�9��9r+9$�?9C$[9��{9W��9Y֤90�9���9Me�9��9&� :��:�X:�X:��:I� :��9�f�9���9.�9Uפ9ۑ�9��{9$[9�?9�+9��9x   